
/*Produced by NSL Core(version=20240424), IP ARCH, Inc. Tue May 21 04:56:15 2024
 Licensed to :EVALUATION USER*/
/*
 DO NOT USE ANY PART OF THIS FILE FOR COMMERCIAL PRODUCTS. 
*/

module add_all ( p_reset , m_clock , sig , start , goal , dig_w , dig_t0 , dig_t1 , dig_t2 , dig_t3 , dig_t4 , dig_t5 , dig_t6 , dig_t7 , dig_t8 , dig_t9 , dig_t10 , dig_t11 , dig_t12 , dig_t13 , dig_t14 , dig_t15 , dig_t16 , dig_t17 , dig_t18 , dig_t19 , dig_t20 , dig_t21 , dig_t22 , dig_t23 , dig_t24 , dig_t25 , dig_t26 , dig_t27 , dig_t28 , dig_t29 , dig_t30 , dig_t31 , dig_t32 , dig_t33 , dig_t34 , dig_t35 , dig_t36 , dig_t37 , dig_t38 , dig_t39 , dig_t40 , dig_t41 , sg_in17 , sg_in18 , sg_in19 , sg_in20 , sg_in21 , sg_in22 , sg_in23 , sg_in24 , sg_in25 , sg_in26 , sg_in27 , sg_in28 , sg_in29 , sg_in30 , sg_in33 , sg_in34 , sg_in35 , sg_in36 , sg_in37 , sg_in38 , sg_in39 , sg_in40 , sg_in41 , sg_in42 , sg_in43 , sg_in44 , sg_in45 , sg_in46 , sg_in49 , sg_in50 , sg_in51 , sg_in52 , sg_in53 , sg_in54 , sg_in55 , sg_in56 , sg_in57 , sg_in58 , sg_in59 , sg_in60 , sg_in61 , sg_in62 , sg_in65 , sg_in66 , sg_in67 , sg_in68 , sg_in69 , sg_in70 , sg_in71 , sg_in72 , sg_in73 , sg_in74 , sg_in75 , sg_in76 , sg_in77 , sg_in78 , sg_in81 , sg_in82 , sg_in83 , sg_in84 , sg_in85 , sg_in86 , sg_in87 , sg_in88 , sg_in89 , sg_in90 , sg_in91 , sg_in92 , sg_in93 , sg_in94 , sg_in97 , sg_in98 , sg_in99 , sg_in100 , sg_in101 , sg_in102 , sg_in103 , sg_in104 , sg_in105 , sg_in106 , sg_in107 , sg_in108 , sg_in109 , sg_in110 , wall_end_in , wall_end , all_sg_in17 , all_sg_in18 , all_sg_in19 , all_sg_in20 , all_sg_in21 , all_sg_in22 , all_sg_in23 , all_sg_in24 , all_sg_in25 , all_sg_in26 , all_sg_in27 , all_sg_in28 , all_sg_in29 , all_sg_in30 , all_sg_in33 , all_sg_in34 , all_sg_in35 , all_sg_in36 , all_sg_in37 , all_sg_in38 , all_sg_in39 , all_sg_in40 , all_sg_in41 , all_sg_in42 , all_sg_in43 , all_sg_in44 , all_sg_in45 , all_sg_in46 , all_sg_in49 , all_sg_in50 , all_sg_in51 , all_sg_in52 , all_sg_in53 , all_sg_in54 , all_sg_in55 , all_sg_in56 , all_sg_in57 , all_sg_in58 , all_sg_in59 , all_sg_in60 , all_sg_in61 , all_sg_in62 , all_sg_in65 , all_sg_in66 , all_sg_in67 , all_sg_in68 , all_sg_in69 , all_sg_in70 , all_sg_in71 , all_sg_in72 , all_sg_in73 , all_sg_in74 , all_sg_in75 , all_sg_in76 , all_sg_in77 , all_sg_in78 , all_sg_in81 , all_sg_in82 , all_sg_in83 , all_sg_in84 , all_sg_in85 , all_sg_in86 , all_sg_in87 , all_sg_in88 , all_sg_in89 , all_sg_in90 , all_sg_in91 , all_sg_in92 , all_sg_in93 , all_sg_in94 , all_sg_in97 , all_sg_in98 , all_sg_in99 , all_sg_in100 , all_sg_in101 , all_sg_in102 , all_sg_in103 , all_sg_in104 , all_sg_in105 , all_sg_in106 , all_sg_in107 , all_sg_in108 , all_sg_in109 , all_sg_in110 , data_in17 , data_in18 , data_in19 , data_in20 , data_in21 , data_in22 , data_in23 , data_in24 , data_in25 , data_in26 , data_in27 , data_in28 , data_in29 , data_in30 , data_in33 , data_in34 , data_in35 , data_in36 , data_in37 , data_in38 , data_in39 , data_in40 , data_in41 , data_in42 , data_in43 , data_in44 , data_in45 , data_in46 , data_in49 , data_in50 , data_in51 , data_in52 , data_in53 , data_in54 , data_in55 , data_in56 , data_in57 , data_in58 , data_in59 , data_in60 , data_in61 , data_in62 , data_in65 , data_in66 , data_in67 , data_in68 , data_in69 , data_in70 , data_in71 , data_in72 , data_in73 , data_in74 , data_in75 , data_in76 , data_in77 , data_in78 , data_in81 , data_in82 , data_in83 , data_in84 , data_in85 , data_in86 , data_in87 , data_in88 , data_in89 , data_in90 , data_in91 , data_in92 , data_in93 , data_in94 , data_in97 , data_in98 , data_in99 , data_in100 , data_in101 , data_in102 , data_in103 , data_in104 , data_in105 , data_in106 , data_in107 , data_in108 , data_in109 , data_in110 , data_in_org17 , data_in_org18 , data_in_org19 , data_in_org20 , data_in_org21 , data_in_org22 , data_in_org23 , data_in_org24 , data_in_org25 , data_in_org26 , data_in_org27 , data_in_org28 , data_in_org29 , data_in_org30 , data_in_org33 , data_in_org34 , data_in_org35 , data_in_org36 , data_in_org37 , data_in_org38 , data_in_org39 , data_in_org40 , data_in_org41 , data_in_org42 , data_in_org43 , data_in_org44 , data_in_org45 , data_in_org46 , data_in_org49 , data_in_org50 , data_in_org51 , data_in_org52 , data_in_org53 , data_in_org54 , data_in_org55 , data_in_org56 , data_in_org57 , data_in_org58 , data_in_org59 , data_in_org60 , data_in_org61 , data_in_org62 , data_in_org65 , data_in_org66 , data_in_org67 , data_in_org68 , data_in_org69 , data_in_org70 , data_in_org71 , data_in_org72 , data_in_org73 , data_in_org74 , data_in_org75 , data_in_org76 , data_in_org77 , data_in_org78 , data_in_org81 , data_in_org82 , data_in_org83 , data_in_org84 , data_in_org85 , data_in_org86 , data_in_org87 , data_in_org88 , data_in_org89 , data_in_org90 , data_in_org91 , data_in_org92 , data_in_org93 , data_in_org94 , data_in_org97 , data_in_org98 , data_in_org99 , data_in_org100 , data_in_org101 , data_in_org102 , data_in_org103 , data_in_org104 , data_in_org105 , data_in_org106 , data_in_org107 , data_in_org108 , data_in_org109 , data_in_org110 , data_out_org17 , data_out_org18 , data_out_org19 , data_out_org20 , data_out_org21 , data_out_org22 , data_out_org23 , data_out_org24 , data_out_org25 , data_out_org26 , data_out_org27 , data_out_org28 , data_out_org29 , data_out_org30 , data_out_org33 , data_out_org34 , data_out_org35 , data_out_org36 , data_out_org37 , data_out_org38 , data_out_org39 , data_out_org40 , data_out_org41 , data_out_org42 , data_out_org43 , data_out_org44 , data_out_org45 , data_out_org46 , data_out_org49 , data_out_org50 , data_out_org51 , data_out_org52 , data_out_org53 , data_out_org54 , data_out_org55 , data_out_org56 , data_out_org57 , data_out_org58 , data_out_org59 , data_out_org60 , data_out_org61 , data_out_org62 , data_out_org65 , data_out_org66 , data_out_org67 , data_out_org68 , data_out_org69 , data_out_org70 , data_out_org71 , data_out_org72 , data_out_org73 , data_out_org74 , data_out_org75 , data_out_org76 , data_out_org77 , data_out_org78 , data_out_org81 , data_out_org82 , data_out_org83 , data_out_org84 , data_out_org85 , data_out_org86 , data_out_org87 , data_out_org88 , data_out_org89 , data_out_org90 , data_out_org91 , data_out_org92 , data_out_org93 , data_out_org94 , data_out_org97 , data_out_org98 , data_out_org99 , data_out_org100 , data_out_org101 , data_out_org102 , data_out_org103 , data_out_org104 , data_out_org105 , data_out_org106 , data_out_org107 , data_out_org108 , data_out_org109 , data_out_org110 , sg_out17 , sg_out18 , sg_out19 , sg_out20 , sg_out21 , sg_out22 , sg_out23 , sg_out24 , sg_out25 , sg_out26 , sg_out27 , sg_out28 , sg_out29 , sg_out30 , sg_out33 , sg_out34 , sg_out35 , sg_out36 , sg_out37 , sg_out38 , sg_out39 , sg_out40 , sg_out41 , sg_out42 , sg_out43 , sg_out44 , sg_out45 , sg_out46 , sg_out49 , sg_out50 , sg_out51 , sg_out52 , sg_out53 , sg_out54 , sg_out55 , sg_out56 , sg_out57 , sg_out58 , sg_out59 , sg_out60 , sg_out61 , sg_out62 , sg_out65 , sg_out66 , sg_out67 , sg_out68 , sg_out69 , sg_out70 , sg_out71 , sg_out72 , sg_out73 , sg_out74 , sg_out75 , sg_out76 , sg_out77 , sg_out78 , sg_out81 , sg_out82 , sg_out83 , sg_out84 , sg_out85 , sg_out86 , sg_out87 , sg_out88 , sg_out89 , sg_out90 , sg_out91 , sg_out92 , sg_out93 , sg_out94 , sg_out97 , sg_out98 , sg_out99 , sg_out100 , sg_out101 , sg_out102 , sg_out103 , sg_out104 , sg_out105 , sg_out106 , sg_out107 , sg_out108 , sg_out109 , sg_out110 , data_out17 , data_out18 , data_out19 , data_out20 , data_out21 , data_out22 , data_out23 , data_out24 , data_out25 , data_out26 , data_out27 , data_out28 , data_out29 , data_out30 , data_out33 , data_out34 , data_out35 , data_out36 , data_out37 , data_out38 , data_out39 , data_out40 , data_out41 , data_out42 , data_out43 , data_out44 , data_out45 , data_out46 , data_out49 , data_out50 , data_out51 , data_out52 , data_out53 , data_out54 , data_out55 , data_out56 , data_out57 , data_out58 , data_out59 , data_out60 , data_out61 , data_out62 , data_out65 , data_out66 , data_out67 , data_out68 , data_out69 , data_out70 , data_out71 , data_out72 , data_out73 , data_out74 , data_out75 , data_out76 , data_out77 , data_out78 , data_out81 , data_out82 , data_out83 , data_out84 , data_out85 , data_out86 , data_out87 , data_out88 , data_out89 , data_out90 , data_out91 , data_out92 , data_out93 , data_out94 , data_out97 , data_out98 , data_out99 , data_out100 , data_out101 , data_out102 , data_out103 , data_out104 , data_out105 , data_out106 , data_out107 , data_out108 , data_out109 , data_out110 , data_out_index17 , data_out_index18 , data_out_index19 , data_out_index20 , data_out_index21 , data_out_index22 , data_out_index23 , data_out_index24 , data_out_index25 , data_out_index26 , data_out_index27 , data_out_index28 , data_out_index29 , data_out_index30 , data_out_index33 , data_out_index34 , data_out_index35 , data_out_index36 , data_out_index37 , data_out_index38 , data_out_index39 , data_out_index40 , data_out_index41 , data_out_index42 , data_out_index43 , data_out_index44 , data_out_index45 , data_out_index46 , data_out_index49 , data_out_index50 , data_out_index51 , data_out_index52 , data_out_index53 , data_out_index54 , data_out_index55 , data_out_index56 , data_out_index57 , data_out_index58 , data_out_index59 , data_out_index60 , data_out_index61 , data_out_index62 , data_out_index65 , data_out_index66 , data_out_index67 , data_out_index68 , data_out_index69 , data_out_index70 , data_out_index71 , data_out_index72 , data_out_index73 , data_out_index74 , data_out_index75 , data_out_index76 , data_out_index77 , data_out_index78 , data_out_index81 , data_out_index82 , data_out_index83 , data_out_index84 , data_out_index85 , data_out_index86 , data_out_index87 , data_out_index88 , data_out_index89 , data_out_index90 , data_out_index91 , data_out_index92 , data_out_index93 , data_out_index94 , data_out_index97 , data_out_index98 , data_out_index99 , data_out_index100 , data_out_index101 , data_out_index102 , data_out_index103 , data_out_index104 , data_out_index105 , data_out_index106 , data_out_index107 , data_out_index108 , data_out_index109 , data_out_index110 , distance_count_all , all_sg_out17 , all_sg_out18 , all_sg_out19 , all_sg_out20 , all_sg_out21 , all_sg_out22 , all_sg_out23 , all_sg_out24 , all_sg_out25 , all_sg_out26 , all_sg_out27 , all_sg_out28 , all_sg_out29 , all_sg_out30 , all_sg_out33 , all_sg_out34 , all_sg_out35 , all_sg_out36 , all_sg_out37 , all_sg_out38 , all_sg_out39 , all_sg_out40 , all_sg_out41 , all_sg_out42 , all_sg_out43 , all_sg_out44 , all_sg_out45 , all_sg_out46 , all_sg_out49 , all_sg_out50 , all_sg_out51 , all_sg_out52 , all_sg_out53 , all_sg_out54 , all_sg_out55 , all_sg_out56 , all_sg_out57 , all_sg_out58 , all_sg_out59 , all_sg_out60 , all_sg_out61 , all_sg_out62 , all_sg_out65 , all_sg_out66 , all_sg_out67 , all_sg_out68 , all_sg_out69 , all_sg_out70 , all_sg_out71 , all_sg_out72 , all_sg_out73 , all_sg_out74 , all_sg_out75 , all_sg_out76 , all_sg_out77 , all_sg_out78 , all_sg_out81 , all_sg_out82 , all_sg_out83 , all_sg_out84 , all_sg_out85 , all_sg_out86 , all_sg_out87 , all_sg_out88 , all_sg_out89 , all_sg_out90 , all_sg_out91 , all_sg_out92 , all_sg_out93 , all_sg_out94 , all_sg_out97 , all_sg_out98 , all_sg_out99 , all_sg_out100 , all_sg_out101 , all_sg_out102 , all_sg_out103 , all_sg_out104 , all_sg_out105 , all_sg_out106 , all_sg_out107 , all_sg_out108 , all_sg_out109 , all_sg_out110 , in_do , out_do , out_data );
  input p_reset, m_clock;
  wire p_reset, m_clock;
  input sig;
  wire sig;
  input [7:0] start;
  wire [7:0] start;
  input [7:0] goal;
  wire [7:0] goal;
  input dig_w;
  wire dig_w;
  output dig_t0;
  wire dig_t0;
  output dig_t1;
  wire dig_t1;
  output dig_t2;
  wire dig_t2;
  output dig_t3;
  wire dig_t3;
  output dig_t4;
  wire dig_t4;
  output dig_t5;
  wire dig_t5;
  output dig_t6;
  wire dig_t6;
  output dig_t7;
  wire dig_t7;
  output dig_t8;
  wire dig_t8;
  output dig_t9;
  wire dig_t9;
  output dig_t10;
  wire dig_t10;
  output dig_t11;
  wire dig_t11;
  output dig_t12;
  wire dig_t12;
  output dig_t13;
  wire dig_t13;
  output dig_t14;
  wire dig_t14;
  output dig_t15;
  wire dig_t15;
  output dig_t16;
  wire dig_t16;
  output dig_t17;
  wire dig_t17;
  output dig_t18;
  wire dig_t18;
  output dig_t19;
  wire dig_t19;
  output dig_t20;
  wire dig_t20;
  output dig_t21;
  wire dig_t21;
  output dig_t22;
  wire dig_t22;
  output dig_t23;
  wire dig_t23;
  output dig_t24;
  wire dig_t24;
  output dig_t25;
  wire dig_t25;
  output dig_t26;
  wire dig_t26;
  output dig_t27;
  wire dig_t27;
  output dig_t28;
  wire dig_t28;
  output dig_t29;
  wire dig_t29;
  output dig_t30;
  wire dig_t30;
  output dig_t31;
  wire dig_t31;
  output dig_t32;
  wire dig_t32;
  output dig_t33;
  wire dig_t33;
  output dig_t34;
  wire dig_t34;
  output dig_t35;
  wire dig_t35;
  output dig_t36;
  wire dig_t36;
  output dig_t37;
  wire dig_t37;
  output dig_t38;
  wire dig_t38;
  output dig_t39;
  wire dig_t39;
  output dig_t40;
  wire dig_t40;
  output dig_t41;
  wire dig_t41;
  input [1:0] sg_in17;
  wire [1:0] sg_in17;
  input [1:0] sg_in18;
  wire [1:0] sg_in18;
  input [1:0] sg_in19;
  wire [1:0] sg_in19;
  input [1:0] sg_in20;
  wire [1:0] sg_in20;
  input [1:0] sg_in21;
  wire [1:0] sg_in21;
  input [1:0] sg_in22;
  wire [1:0] sg_in22;
  input [1:0] sg_in23;
  wire [1:0] sg_in23;
  input [1:0] sg_in24;
  wire [1:0] sg_in24;
  input [1:0] sg_in25;
  wire [1:0] sg_in25;
  input [1:0] sg_in26;
  wire [1:0] sg_in26;
  input [1:0] sg_in27;
  wire [1:0] sg_in27;
  input [1:0] sg_in28;
  wire [1:0] sg_in28;
  input [1:0] sg_in29;
  wire [1:0] sg_in29;
  input [1:0] sg_in30;
  wire [1:0] sg_in30;
  input [1:0] sg_in33;
  wire [1:0] sg_in33;
  input [1:0] sg_in34;
  wire [1:0] sg_in34;
  input [1:0] sg_in35;
  wire [1:0] sg_in35;
  input [1:0] sg_in36;
  wire [1:0] sg_in36;
  input [1:0] sg_in37;
  wire [1:0] sg_in37;
  input [1:0] sg_in38;
  wire [1:0] sg_in38;
  input [1:0] sg_in39;
  wire [1:0] sg_in39;
  input [1:0] sg_in40;
  wire [1:0] sg_in40;
  input [1:0] sg_in41;
  wire [1:0] sg_in41;
  input [1:0] sg_in42;
  wire [1:0] sg_in42;
  input [1:0] sg_in43;
  wire [1:0] sg_in43;
  input [1:0] sg_in44;
  wire [1:0] sg_in44;
  input [1:0] sg_in45;
  wire [1:0] sg_in45;
  input [1:0] sg_in46;
  wire [1:0] sg_in46;
  input [1:0] sg_in49;
  wire [1:0] sg_in49;
  input [1:0] sg_in50;
  wire [1:0] sg_in50;
  input [1:0] sg_in51;
  wire [1:0] sg_in51;
  input [1:0] sg_in52;
  wire [1:0] sg_in52;
  input [1:0] sg_in53;
  wire [1:0] sg_in53;
  input [1:0] sg_in54;
  wire [1:0] sg_in54;
  input [1:0] sg_in55;
  wire [1:0] sg_in55;
  input [1:0] sg_in56;
  wire [1:0] sg_in56;
  input [1:0] sg_in57;
  wire [1:0] sg_in57;
  input [1:0] sg_in58;
  wire [1:0] sg_in58;
  input [1:0] sg_in59;
  wire [1:0] sg_in59;
  input [1:0] sg_in60;
  wire [1:0] sg_in60;
  input [1:0] sg_in61;
  wire [1:0] sg_in61;
  input [1:0] sg_in62;
  wire [1:0] sg_in62;
  input [1:0] sg_in65;
  wire [1:0] sg_in65;
  input [1:0] sg_in66;
  wire [1:0] sg_in66;
  input [1:0] sg_in67;
  wire [1:0] sg_in67;
  input [1:0] sg_in68;
  wire [1:0] sg_in68;
  input [1:0] sg_in69;
  wire [1:0] sg_in69;
  input [1:0] sg_in70;
  wire [1:0] sg_in70;
  input [1:0] sg_in71;
  wire [1:0] sg_in71;
  input [1:0] sg_in72;
  wire [1:0] sg_in72;
  input [1:0] sg_in73;
  wire [1:0] sg_in73;
  input [1:0] sg_in74;
  wire [1:0] sg_in74;
  input [1:0] sg_in75;
  wire [1:0] sg_in75;
  input [1:0] sg_in76;
  wire [1:0] sg_in76;
  input [1:0] sg_in77;
  wire [1:0] sg_in77;
  input [1:0] sg_in78;
  wire [1:0] sg_in78;
  input [1:0] sg_in81;
  wire [1:0] sg_in81;
  input [1:0] sg_in82;
  wire [1:0] sg_in82;
  input [1:0] sg_in83;
  wire [1:0] sg_in83;
  input [1:0] sg_in84;
  wire [1:0] sg_in84;
  input [1:0] sg_in85;
  wire [1:0] sg_in85;
  input [1:0] sg_in86;
  wire [1:0] sg_in86;
  input [1:0] sg_in87;
  wire [1:0] sg_in87;
  input [1:0] sg_in88;
  wire [1:0] sg_in88;
  input [1:0] sg_in89;
  wire [1:0] sg_in89;
  input [1:0] sg_in90;
  wire [1:0] sg_in90;
  input [1:0] sg_in91;
  wire [1:0] sg_in91;
  input [1:0] sg_in92;
  wire [1:0] sg_in92;
  input [1:0] sg_in93;
  wire [1:0] sg_in93;
  input [1:0] sg_in94;
  wire [1:0] sg_in94;
  input [1:0] sg_in97;
  wire [1:0] sg_in97;
  input [1:0] sg_in98;
  wire [1:0] sg_in98;
  input [1:0] sg_in99;
  wire [1:0] sg_in99;
  input [1:0] sg_in100;
  wire [1:0] sg_in100;
  input [1:0] sg_in101;
  wire [1:0] sg_in101;
  input [1:0] sg_in102;
  wire [1:0] sg_in102;
  input [1:0] sg_in103;
  wire [1:0] sg_in103;
  input [1:0] sg_in104;
  wire [1:0] sg_in104;
  input [1:0] sg_in105;
  wire [1:0] sg_in105;
  input [1:0] sg_in106;
  wire [1:0] sg_in106;
  input [1:0] sg_in107;
  wire [1:0] sg_in107;
  input [1:0] sg_in108;
  wire [1:0] sg_in108;
  input [1:0] sg_in109;
  wire [1:0] sg_in109;
  input [1:0] sg_in110;
  wire [1:0] sg_in110;
  input [127:0] wall_end_in;
  wire [127:0] wall_end_in;
  output [127:0] wall_end;
  wire [127:0] wall_end;
  input [127:0] all_sg_in17;
  wire [127:0] all_sg_in17;
  input [127:0] all_sg_in18;
  wire [127:0] all_sg_in18;
  input [127:0] all_sg_in19;
  wire [127:0] all_sg_in19;
  input [127:0] all_sg_in20;
  wire [127:0] all_sg_in20;
  input [127:0] all_sg_in21;
  wire [127:0] all_sg_in21;
  input [127:0] all_sg_in22;
  wire [127:0] all_sg_in22;
  input [127:0] all_sg_in23;
  wire [127:0] all_sg_in23;
  input [127:0] all_sg_in24;
  wire [127:0] all_sg_in24;
  input [127:0] all_sg_in25;
  wire [127:0] all_sg_in25;
  input [127:0] all_sg_in26;
  wire [127:0] all_sg_in26;
  input [127:0] all_sg_in27;
  wire [127:0] all_sg_in27;
  input [127:0] all_sg_in28;
  wire [127:0] all_sg_in28;
  input [127:0] all_sg_in29;
  wire [127:0] all_sg_in29;
  input [127:0] all_sg_in30;
  wire [127:0] all_sg_in30;
  input [127:0] all_sg_in33;
  wire [127:0] all_sg_in33;
  input [127:0] all_sg_in34;
  wire [127:0] all_sg_in34;
  input [127:0] all_sg_in35;
  wire [127:0] all_sg_in35;
  input [127:0] all_sg_in36;
  wire [127:0] all_sg_in36;
  input [127:0] all_sg_in37;
  wire [127:0] all_sg_in37;
  input [127:0] all_sg_in38;
  wire [127:0] all_sg_in38;
  input [127:0] all_sg_in39;
  wire [127:0] all_sg_in39;
  input [127:0] all_sg_in40;
  wire [127:0] all_sg_in40;
  input [127:0] all_sg_in41;
  wire [127:0] all_sg_in41;
  input [127:0] all_sg_in42;
  wire [127:0] all_sg_in42;
  input [127:0] all_sg_in43;
  wire [127:0] all_sg_in43;
  input [127:0] all_sg_in44;
  wire [127:0] all_sg_in44;
  input [127:0] all_sg_in45;
  wire [127:0] all_sg_in45;
  input [127:0] all_sg_in46;
  wire [127:0] all_sg_in46;
  input [127:0] all_sg_in49;
  wire [127:0] all_sg_in49;
  input [127:0] all_sg_in50;
  wire [127:0] all_sg_in50;
  input [127:0] all_sg_in51;
  wire [127:0] all_sg_in51;
  input [127:0] all_sg_in52;
  wire [127:0] all_sg_in52;
  input [127:0] all_sg_in53;
  wire [127:0] all_sg_in53;
  input [127:0] all_sg_in54;
  wire [127:0] all_sg_in54;
  input [127:0] all_sg_in55;
  wire [127:0] all_sg_in55;
  input [127:0] all_sg_in56;
  wire [127:0] all_sg_in56;
  input [127:0] all_sg_in57;
  wire [127:0] all_sg_in57;
  input [127:0] all_sg_in58;
  wire [127:0] all_sg_in58;
  input [127:0] all_sg_in59;
  wire [127:0] all_sg_in59;
  input [127:0] all_sg_in60;
  wire [127:0] all_sg_in60;
  input [127:0] all_sg_in61;
  wire [127:0] all_sg_in61;
  input [127:0] all_sg_in62;
  wire [127:0] all_sg_in62;
  input [127:0] all_sg_in65;
  wire [127:0] all_sg_in65;
  input [127:0] all_sg_in66;
  wire [127:0] all_sg_in66;
  input [127:0] all_sg_in67;
  wire [127:0] all_sg_in67;
  input [127:0] all_sg_in68;
  wire [127:0] all_sg_in68;
  input [127:0] all_sg_in69;
  wire [127:0] all_sg_in69;
  input [127:0] all_sg_in70;
  wire [127:0] all_sg_in70;
  input [127:0] all_sg_in71;
  wire [127:0] all_sg_in71;
  input [127:0] all_sg_in72;
  wire [127:0] all_sg_in72;
  input [127:0] all_sg_in73;
  wire [127:0] all_sg_in73;
  input [127:0] all_sg_in74;
  wire [127:0] all_sg_in74;
  input [127:0] all_sg_in75;
  wire [127:0] all_sg_in75;
  input [127:0] all_sg_in76;
  wire [127:0] all_sg_in76;
  input [127:0] all_sg_in77;
  wire [127:0] all_sg_in77;
  input [127:0] all_sg_in78;
  wire [127:0] all_sg_in78;
  input [127:0] all_sg_in81;
  wire [127:0] all_sg_in81;
  input [127:0] all_sg_in82;
  wire [127:0] all_sg_in82;
  input [127:0] all_sg_in83;
  wire [127:0] all_sg_in83;
  input [127:0] all_sg_in84;
  wire [127:0] all_sg_in84;
  input [127:0] all_sg_in85;
  wire [127:0] all_sg_in85;
  input [127:0] all_sg_in86;
  wire [127:0] all_sg_in86;
  input [127:0] all_sg_in87;
  wire [127:0] all_sg_in87;
  input [127:0] all_sg_in88;
  wire [127:0] all_sg_in88;
  input [127:0] all_sg_in89;
  wire [127:0] all_sg_in89;
  input [127:0] all_sg_in90;
  wire [127:0] all_sg_in90;
  input [127:0] all_sg_in91;
  wire [127:0] all_sg_in91;
  input [127:0] all_sg_in92;
  wire [127:0] all_sg_in92;
  input [127:0] all_sg_in93;
  wire [127:0] all_sg_in93;
  input [127:0] all_sg_in94;
  wire [127:0] all_sg_in94;
  input [127:0] all_sg_in97;
  wire [127:0] all_sg_in97;
  input [127:0] all_sg_in98;
  wire [127:0] all_sg_in98;
  input [127:0] all_sg_in99;
  wire [127:0] all_sg_in99;
  input [127:0] all_sg_in100;
  wire [127:0] all_sg_in100;
  input [127:0] all_sg_in101;
  wire [127:0] all_sg_in101;
  input [127:0] all_sg_in102;
  wire [127:0] all_sg_in102;
  input [127:0] all_sg_in103;
  wire [127:0] all_sg_in103;
  input [127:0] all_sg_in104;
  wire [127:0] all_sg_in104;
  input [127:0] all_sg_in105;
  wire [127:0] all_sg_in105;
  input [127:0] all_sg_in106;
  wire [127:0] all_sg_in106;
  input [127:0] all_sg_in107;
  wire [127:0] all_sg_in107;
  input [127:0] all_sg_in108;
  wire [127:0] all_sg_in108;
  input [127:0] all_sg_in109;
  wire [127:0] all_sg_in109;
  input [127:0] all_sg_in110;
  wire [127:0] all_sg_in110;
  input [7:0] data_in17;
  wire [7:0] data_in17;
  input [7:0] data_in18;
  wire [7:0] data_in18;
  input [7:0] data_in19;
  wire [7:0] data_in19;
  input [7:0] data_in20;
  wire [7:0] data_in20;
  input [7:0] data_in21;
  wire [7:0] data_in21;
  input [7:0] data_in22;
  wire [7:0] data_in22;
  input [7:0] data_in23;
  wire [7:0] data_in23;
  input [7:0] data_in24;
  wire [7:0] data_in24;
  input [7:0] data_in25;
  wire [7:0] data_in25;
  input [7:0] data_in26;
  wire [7:0] data_in26;
  input [7:0] data_in27;
  wire [7:0] data_in27;
  input [7:0] data_in28;
  wire [7:0] data_in28;
  input [7:0] data_in29;
  wire [7:0] data_in29;
  input [7:0] data_in30;
  wire [7:0] data_in30;
  input [7:0] data_in33;
  wire [7:0] data_in33;
  input [7:0] data_in34;
  wire [7:0] data_in34;
  input [7:0] data_in35;
  wire [7:0] data_in35;
  input [7:0] data_in36;
  wire [7:0] data_in36;
  input [7:0] data_in37;
  wire [7:0] data_in37;
  input [7:0] data_in38;
  wire [7:0] data_in38;
  input [7:0] data_in39;
  wire [7:0] data_in39;
  input [7:0] data_in40;
  wire [7:0] data_in40;
  input [7:0] data_in41;
  wire [7:0] data_in41;
  input [7:0] data_in42;
  wire [7:0] data_in42;
  input [7:0] data_in43;
  wire [7:0] data_in43;
  input [7:0] data_in44;
  wire [7:0] data_in44;
  input [7:0] data_in45;
  wire [7:0] data_in45;
  input [7:0] data_in46;
  wire [7:0] data_in46;
  input [7:0] data_in49;
  wire [7:0] data_in49;
  input [7:0] data_in50;
  wire [7:0] data_in50;
  input [7:0] data_in51;
  wire [7:0] data_in51;
  input [7:0] data_in52;
  wire [7:0] data_in52;
  input [7:0] data_in53;
  wire [7:0] data_in53;
  input [7:0] data_in54;
  wire [7:0] data_in54;
  input [7:0] data_in55;
  wire [7:0] data_in55;
  input [7:0] data_in56;
  wire [7:0] data_in56;
  input [7:0] data_in57;
  wire [7:0] data_in57;
  input [7:0] data_in58;
  wire [7:0] data_in58;
  input [7:0] data_in59;
  wire [7:0] data_in59;
  input [7:0] data_in60;
  wire [7:0] data_in60;
  input [7:0] data_in61;
  wire [7:0] data_in61;
  input [7:0] data_in62;
  wire [7:0] data_in62;
  input [7:0] data_in65;
  wire [7:0] data_in65;
  input [7:0] data_in66;
  wire [7:0] data_in66;
  input [7:0] data_in67;
  wire [7:0] data_in67;
  input [7:0] data_in68;
  wire [7:0] data_in68;
  input [7:0] data_in69;
  wire [7:0] data_in69;
  input [7:0] data_in70;
  wire [7:0] data_in70;
  input [7:0] data_in71;
  wire [7:0] data_in71;
  input [7:0] data_in72;
  wire [7:0] data_in72;
  input [7:0] data_in73;
  wire [7:0] data_in73;
  input [7:0] data_in74;
  wire [7:0] data_in74;
  input [7:0] data_in75;
  wire [7:0] data_in75;
  input [7:0] data_in76;
  wire [7:0] data_in76;
  input [7:0] data_in77;
  wire [7:0] data_in77;
  input [7:0] data_in78;
  wire [7:0] data_in78;
  input [7:0] data_in81;
  wire [7:0] data_in81;
  input [7:0] data_in82;
  wire [7:0] data_in82;
  input [7:0] data_in83;
  wire [7:0] data_in83;
  input [7:0] data_in84;
  wire [7:0] data_in84;
  input [7:0] data_in85;
  wire [7:0] data_in85;
  input [7:0] data_in86;
  wire [7:0] data_in86;
  input [7:0] data_in87;
  wire [7:0] data_in87;
  input [7:0] data_in88;
  wire [7:0] data_in88;
  input [7:0] data_in89;
  wire [7:0] data_in89;
  input [7:0] data_in90;
  wire [7:0] data_in90;
  input [7:0] data_in91;
  wire [7:0] data_in91;
  input [7:0] data_in92;
  wire [7:0] data_in92;
  input [7:0] data_in93;
  wire [7:0] data_in93;
  input [7:0] data_in94;
  wire [7:0] data_in94;
  input [7:0] data_in97;
  wire [7:0] data_in97;
  input [7:0] data_in98;
  wire [7:0] data_in98;
  input [7:0] data_in99;
  wire [7:0] data_in99;
  input [7:0] data_in100;
  wire [7:0] data_in100;
  input [7:0] data_in101;
  wire [7:0] data_in101;
  input [7:0] data_in102;
  wire [7:0] data_in102;
  input [7:0] data_in103;
  wire [7:0] data_in103;
  input [7:0] data_in104;
  wire [7:0] data_in104;
  input [7:0] data_in105;
  wire [7:0] data_in105;
  input [7:0] data_in106;
  wire [7:0] data_in106;
  input [7:0] data_in107;
  wire [7:0] data_in107;
  input [7:0] data_in108;
  wire [7:0] data_in108;
  input [7:0] data_in109;
  wire [7:0] data_in109;
  input [7:0] data_in110;
  wire [7:0] data_in110;
  input [7:0] data_in_org17;
  wire [7:0] data_in_org17;
  input [7:0] data_in_org18;
  wire [7:0] data_in_org18;
  input [7:0] data_in_org19;
  wire [7:0] data_in_org19;
  input [7:0] data_in_org20;
  wire [7:0] data_in_org20;
  input [7:0] data_in_org21;
  wire [7:0] data_in_org21;
  input [7:0] data_in_org22;
  wire [7:0] data_in_org22;
  input [7:0] data_in_org23;
  wire [7:0] data_in_org23;
  input [7:0] data_in_org24;
  wire [7:0] data_in_org24;
  input [7:0] data_in_org25;
  wire [7:0] data_in_org25;
  input [7:0] data_in_org26;
  wire [7:0] data_in_org26;
  input [7:0] data_in_org27;
  wire [7:0] data_in_org27;
  input [7:0] data_in_org28;
  wire [7:0] data_in_org28;
  input [7:0] data_in_org29;
  wire [7:0] data_in_org29;
  input [7:0] data_in_org30;
  wire [7:0] data_in_org30;
  input [7:0] data_in_org33;
  wire [7:0] data_in_org33;
  input [7:0] data_in_org34;
  wire [7:0] data_in_org34;
  input [7:0] data_in_org35;
  wire [7:0] data_in_org35;
  input [7:0] data_in_org36;
  wire [7:0] data_in_org36;
  input [7:0] data_in_org37;
  wire [7:0] data_in_org37;
  input [7:0] data_in_org38;
  wire [7:0] data_in_org38;
  input [7:0] data_in_org39;
  wire [7:0] data_in_org39;
  input [7:0] data_in_org40;
  wire [7:0] data_in_org40;
  input [7:0] data_in_org41;
  wire [7:0] data_in_org41;
  input [7:0] data_in_org42;
  wire [7:0] data_in_org42;
  input [7:0] data_in_org43;
  wire [7:0] data_in_org43;
  input [7:0] data_in_org44;
  wire [7:0] data_in_org44;
  input [7:0] data_in_org45;
  wire [7:0] data_in_org45;
  input [7:0] data_in_org46;
  wire [7:0] data_in_org46;
  input [7:0] data_in_org49;
  wire [7:0] data_in_org49;
  input [7:0] data_in_org50;
  wire [7:0] data_in_org50;
  input [7:0] data_in_org51;
  wire [7:0] data_in_org51;
  input [7:0] data_in_org52;
  wire [7:0] data_in_org52;
  input [7:0] data_in_org53;
  wire [7:0] data_in_org53;
  input [7:0] data_in_org54;
  wire [7:0] data_in_org54;
  input [7:0] data_in_org55;
  wire [7:0] data_in_org55;
  input [7:0] data_in_org56;
  wire [7:0] data_in_org56;
  input [7:0] data_in_org57;
  wire [7:0] data_in_org57;
  input [7:0] data_in_org58;
  wire [7:0] data_in_org58;
  input [7:0] data_in_org59;
  wire [7:0] data_in_org59;
  input [7:0] data_in_org60;
  wire [7:0] data_in_org60;
  input [7:0] data_in_org61;
  wire [7:0] data_in_org61;
  input [7:0] data_in_org62;
  wire [7:0] data_in_org62;
  input [7:0] data_in_org65;
  wire [7:0] data_in_org65;
  input [7:0] data_in_org66;
  wire [7:0] data_in_org66;
  input [7:0] data_in_org67;
  wire [7:0] data_in_org67;
  input [7:0] data_in_org68;
  wire [7:0] data_in_org68;
  input [7:0] data_in_org69;
  wire [7:0] data_in_org69;
  input [7:0] data_in_org70;
  wire [7:0] data_in_org70;
  input [7:0] data_in_org71;
  wire [7:0] data_in_org71;
  input [7:0] data_in_org72;
  wire [7:0] data_in_org72;
  input [7:0] data_in_org73;
  wire [7:0] data_in_org73;
  input [7:0] data_in_org74;
  wire [7:0] data_in_org74;
  input [7:0] data_in_org75;
  wire [7:0] data_in_org75;
  input [7:0] data_in_org76;
  wire [7:0] data_in_org76;
  input [7:0] data_in_org77;
  wire [7:0] data_in_org77;
  input [7:0] data_in_org78;
  wire [7:0] data_in_org78;
  input [7:0] data_in_org81;
  wire [7:0] data_in_org81;
  input [7:0] data_in_org82;
  wire [7:0] data_in_org82;
  input [7:0] data_in_org83;
  wire [7:0] data_in_org83;
  input [7:0] data_in_org84;
  wire [7:0] data_in_org84;
  input [7:0] data_in_org85;
  wire [7:0] data_in_org85;
  input [7:0] data_in_org86;
  wire [7:0] data_in_org86;
  input [7:0] data_in_org87;
  wire [7:0] data_in_org87;
  input [7:0] data_in_org88;
  wire [7:0] data_in_org88;
  input [7:0] data_in_org89;
  wire [7:0] data_in_org89;
  input [7:0] data_in_org90;
  wire [7:0] data_in_org90;
  input [7:0] data_in_org91;
  wire [7:0] data_in_org91;
  input [7:0] data_in_org92;
  wire [7:0] data_in_org92;
  input [7:0] data_in_org93;
  wire [7:0] data_in_org93;
  input [7:0] data_in_org94;
  wire [7:0] data_in_org94;
  input [7:0] data_in_org97;
  wire [7:0] data_in_org97;
  input [7:0] data_in_org98;
  wire [7:0] data_in_org98;
  input [7:0] data_in_org99;
  wire [7:0] data_in_org99;
  input [7:0] data_in_org100;
  wire [7:0] data_in_org100;
  input [7:0] data_in_org101;
  wire [7:0] data_in_org101;
  input [7:0] data_in_org102;
  wire [7:0] data_in_org102;
  input [7:0] data_in_org103;
  wire [7:0] data_in_org103;
  input [7:0] data_in_org104;
  wire [7:0] data_in_org104;
  input [7:0] data_in_org105;
  wire [7:0] data_in_org105;
  input [7:0] data_in_org106;
  wire [7:0] data_in_org106;
  input [7:0] data_in_org107;
  wire [7:0] data_in_org107;
  input [7:0] data_in_org108;
  wire [7:0] data_in_org108;
  input [7:0] data_in_org109;
  wire [7:0] data_in_org109;
  input [7:0] data_in_org110;
  wire [7:0] data_in_org110;
  output [7:0] data_out_org17;
  wire [7:0] data_out_org17;
  output [7:0] data_out_org18;
  wire [7:0] data_out_org18;
  output [7:0] data_out_org19;
  wire [7:0] data_out_org19;
  output [7:0] data_out_org20;
  wire [7:0] data_out_org20;
  output [7:0] data_out_org21;
  wire [7:0] data_out_org21;
  output [7:0] data_out_org22;
  wire [7:0] data_out_org22;
  output [7:0] data_out_org23;
  wire [7:0] data_out_org23;
  output [7:0] data_out_org24;
  wire [7:0] data_out_org24;
  output [7:0] data_out_org25;
  wire [7:0] data_out_org25;
  output [7:0] data_out_org26;
  wire [7:0] data_out_org26;
  output [7:0] data_out_org27;
  wire [7:0] data_out_org27;
  output [7:0] data_out_org28;
  wire [7:0] data_out_org28;
  output [7:0] data_out_org29;
  wire [7:0] data_out_org29;
  output [7:0] data_out_org30;
  wire [7:0] data_out_org30;
  output [7:0] data_out_org33;
  wire [7:0] data_out_org33;
  output [7:0] data_out_org34;
  wire [7:0] data_out_org34;
  output [7:0] data_out_org35;
  wire [7:0] data_out_org35;
  output [7:0] data_out_org36;
  wire [7:0] data_out_org36;
  output [7:0] data_out_org37;
  wire [7:0] data_out_org37;
  output [7:0] data_out_org38;
  wire [7:0] data_out_org38;
  output [7:0] data_out_org39;
  wire [7:0] data_out_org39;
  output [7:0] data_out_org40;
  wire [7:0] data_out_org40;
  output [7:0] data_out_org41;
  wire [7:0] data_out_org41;
  output [7:0] data_out_org42;
  wire [7:0] data_out_org42;
  output [7:0] data_out_org43;
  wire [7:0] data_out_org43;
  output [7:0] data_out_org44;
  wire [7:0] data_out_org44;
  output [7:0] data_out_org45;
  wire [7:0] data_out_org45;
  output [7:0] data_out_org46;
  wire [7:0] data_out_org46;
  output [7:0] data_out_org49;
  wire [7:0] data_out_org49;
  output [7:0] data_out_org50;
  wire [7:0] data_out_org50;
  output [7:0] data_out_org51;
  wire [7:0] data_out_org51;
  output [7:0] data_out_org52;
  wire [7:0] data_out_org52;
  output [7:0] data_out_org53;
  wire [7:0] data_out_org53;
  output [7:0] data_out_org54;
  wire [7:0] data_out_org54;
  output [7:0] data_out_org55;
  wire [7:0] data_out_org55;
  output [7:0] data_out_org56;
  wire [7:0] data_out_org56;
  output [7:0] data_out_org57;
  wire [7:0] data_out_org57;
  output [7:0] data_out_org58;
  wire [7:0] data_out_org58;
  output [7:0] data_out_org59;
  wire [7:0] data_out_org59;
  output [7:0] data_out_org60;
  wire [7:0] data_out_org60;
  output [7:0] data_out_org61;
  wire [7:0] data_out_org61;
  output [7:0] data_out_org62;
  wire [7:0] data_out_org62;
  output [7:0] data_out_org65;
  wire [7:0] data_out_org65;
  output [7:0] data_out_org66;
  wire [7:0] data_out_org66;
  output [7:0] data_out_org67;
  wire [7:0] data_out_org67;
  output [7:0] data_out_org68;
  wire [7:0] data_out_org68;
  output [7:0] data_out_org69;
  wire [7:0] data_out_org69;
  output [7:0] data_out_org70;
  wire [7:0] data_out_org70;
  output [7:0] data_out_org71;
  wire [7:0] data_out_org71;
  output [7:0] data_out_org72;
  wire [7:0] data_out_org72;
  output [7:0] data_out_org73;
  wire [7:0] data_out_org73;
  output [7:0] data_out_org74;
  wire [7:0] data_out_org74;
  output [7:0] data_out_org75;
  wire [7:0] data_out_org75;
  output [7:0] data_out_org76;
  wire [7:0] data_out_org76;
  output [7:0] data_out_org77;
  wire [7:0] data_out_org77;
  output [7:0] data_out_org78;
  wire [7:0] data_out_org78;
  output [7:0] data_out_org81;
  wire [7:0] data_out_org81;
  output [7:0] data_out_org82;
  wire [7:0] data_out_org82;
  output [7:0] data_out_org83;
  wire [7:0] data_out_org83;
  output [7:0] data_out_org84;
  wire [7:0] data_out_org84;
  output [7:0] data_out_org85;
  wire [7:0] data_out_org85;
  output [7:0] data_out_org86;
  wire [7:0] data_out_org86;
  output [7:0] data_out_org87;
  wire [7:0] data_out_org87;
  output [7:0] data_out_org88;
  wire [7:0] data_out_org88;
  output [7:0] data_out_org89;
  wire [7:0] data_out_org89;
  output [7:0] data_out_org90;
  wire [7:0] data_out_org90;
  output [7:0] data_out_org91;
  wire [7:0] data_out_org91;
  output [7:0] data_out_org92;
  wire [7:0] data_out_org92;
  output [7:0] data_out_org93;
  wire [7:0] data_out_org93;
  output [7:0] data_out_org94;
  wire [7:0] data_out_org94;
  output [7:0] data_out_org97;
  wire [7:0] data_out_org97;
  output [7:0] data_out_org98;
  wire [7:0] data_out_org98;
  output [7:0] data_out_org99;
  wire [7:0] data_out_org99;
  output [7:0] data_out_org100;
  wire [7:0] data_out_org100;
  output [7:0] data_out_org101;
  wire [7:0] data_out_org101;
  output [7:0] data_out_org102;
  wire [7:0] data_out_org102;
  output [7:0] data_out_org103;
  wire [7:0] data_out_org103;
  output [7:0] data_out_org104;
  wire [7:0] data_out_org104;
  output [7:0] data_out_org105;
  wire [7:0] data_out_org105;
  output [7:0] data_out_org106;
  wire [7:0] data_out_org106;
  output [7:0] data_out_org107;
  wire [7:0] data_out_org107;
  output [7:0] data_out_org108;
  wire [7:0] data_out_org108;
  output [7:0] data_out_org109;
  wire [7:0] data_out_org109;
  output [7:0] data_out_org110;
  wire [7:0] data_out_org110;
  output [1:0] sg_out17;
  wire [1:0] sg_out17;
  output [1:0] sg_out18;
  wire [1:0] sg_out18;
  output [1:0] sg_out19;
  wire [1:0] sg_out19;
  output [1:0] sg_out20;
  wire [1:0] sg_out20;
  output [1:0] sg_out21;
  wire [1:0] sg_out21;
  output [1:0] sg_out22;
  wire [1:0] sg_out22;
  output [1:0] sg_out23;
  wire [1:0] sg_out23;
  output [1:0] sg_out24;
  wire [1:0] sg_out24;
  output [1:0] sg_out25;
  wire [1:0] sg_out25;
  output [1:0] sg_out26;
  wire [1:0] sg_out26;
  output [1:0] sg_out27;
  wire [1:0] sg_out27;
  output [1:0] sg_out28;
  wire [1:0] sg_out28;
  output [1:0] sg_out29;
  wire [1:0] sg_out29;
  output [1:0] sg_out30;
  wire [1:0] sg_out30;
  output [1:0] sg_out33;
  wire [1:0] sg_out33;
  output [1:0] sg_out34;
  wire [1:0] sg_out34;
  output [1:0] sg_out35;
  wire [1:0] sg_out35;
  output [1:0] sg_out36;
  wire [1:0] sg_out36;
  output [1:0] sg_out37;
  wire [1:0] sg_out37;
  output [1:0] sg_out38;
  wire [1:0] sg_out38;
  output [1:0] sg_out39;
  wire [1:0] sg_out39;
  output [1:0] sg_out40;
  wire [1:0] sg_out40;
  output [1:0] sg_out41;
  wire [1:0] sg_out41;
  output [1:0] sg_out42;
  wire [1:0] sg_out42;
  output [1:0] sg_out43;
  wire [1:0] sg_out43;
  output [1:0] sg_out44;
  wire [1:0] sg_out44;
  output [1:0] sg_out45;
  wire [1:0] sg_out45;
  output [1:0] sg_out46;
  wire [1:0] sg_out46;
  output [1:0] sg_out49;
  wire [1:0] sg_out49;
  output [1:0] sg_out50;
  wire [1:0] sg_out50;
  output [1:0] sg_out51;
  wire [1:0] sg_out51;
  output [1:0] sg_out52;
  wire [1:0] sg_out52;
  output [1:0] sg_out53;
  wire [1:0] sg_out53;
  output [1:0] sg_out54;
  wire [1:0] sg_out54;
  output [1:0] sg_out55;
  wire [1:0] sg_out55;
  output [1:0] sg_out56;
  wire [1:0] sg_out56;
  output [1:0] sg_out57;
  wire [1:0] sg_out57;
  output [1:0] sg_out58;
  wire [1:0] sg_out58;
  output [1:0] sg_out59;
  wire [1:0] sg_out59;
  output [1:0] sg_out60;
  wire [1:0] sg_out60;
  output [1:0] sg_out61;
  wire [1:0] sg_out61;
  output [1:0] sg_out62;
  wire [1:0] sg_out62;
  output [1:0] sg_out65;
  wire [1:0] sg_out65;
  output [1:0] sg_out66;
  wire [1:0] sg_out66;
  output [1:0] sg_out67;
  wire [1:0] sg_out67;
  output [1:0] sg_out68;
  wire [1:0] sg_out68;
  output [1:0] sg_out69;
  wire [1:0] sg_out69;
  output [1:0] sg_out70;
  wire [1:0] sg_out70;
  output [1:0] sg_out71;
  wire [1:0] sg_out71;
  output [1:0] sg_out72;
  wire [1:0] sg_out72;
  output [1:0] sg_out73;
  wire [1:0] sg_out73;
  output [1:0] sg_out74;
  wire [1:0] sg_out74;
  output [1:0] sg_out75;
  wire [1:0] sg_out75;
  output [1:0] sg_out76;
  wire [1:0] sg_out76;
  output [1:0] sg_out77;
  wire [1:0] sg_out77;
  output [1:0] sg_out78;
  wire [1:0] sg_out78;
  output [1:0] sg_out81;
  wire [1:0] sg_out81;
  output [1:0] sg_out82;
  wire [1:0] sg_out82;
  output [1:0] sg_out83;
  wire [1:0] sg_out83;
  output [1:0] sg_out84;
  wire [1:0] sg_out84;
  output [1:0] sg_out85;
  wire [1:0] sg_out85;
  output [1:0] sg_out86;
  wire [1:0] sg_out86;
  output [1:0] sg_out87;
  wire [1:0] sg_out87;
  output [1:0] sg_out88;
  wire [1:0] sg_out88;
  output [1:0] sg_out89;
  wire [1:0] sg_out89;
  output [1:0] sg_out90;
  wire [1:0] sg_out90;
  output [1:0] sg_out91;
  wire [1:0] sg_out91;
  output [1:0] sg_out92;
  wire [1:0] sg_out92;
  output [1:0] sg_out93;
  wire [1:0] sg_out93;
  output [1:0] sg_out94;
  wire [1:0] sg_out94;
  output [1:0] sg_out97;
  wire [1:0] sg_out97;
  output [1:0] sg_out98;
  wire [1:0] sg_out98;
  output [1:0] sg_out99;
  wire [1:0] sg_out99;
  output [1:0] sg_out100;
  wire [1:0] sg_out100;
  output [1:0] sg_out101;
  wire [1:0] sg_out101;
  output [1:0] sg_out102;
  wire [1:0] sg_out102;
  output [1:0] sg_out103;
  wire [1:0] sg_out103;
  output [1:0] sg_out104;
  wire [1:0] sg_out104;
  output [1:0] sg_out105;
  wire [1:0] sg_out105;
  output [1:0] sg_out106;
  wire [1:0] sg_out106;
  output [1:0] sg_out107;
  wire [1:0] sg_out107;
  output [1:0] sg_out108;
  wire [1:0] sg_out108;
  output [1:0] sg_out109;
  wire [1:0] sg_out109;
  output [1:0] sg_out110;
  wire [1:0] sg_out110;
  output [7:0] data_out17;
  wire [7:0] data_out17;
  output [7:0] data_out18;
  wire [7:0] data_out18;
  output [7:0] data_out19;
  wire [7:0] data_out19;
  output [7:0] data_out20;
  wire [7:0] data_out20;
  output [7:0] data_out21;
  wire [7:0] data_out21;
  output [7:0] data_out22;
  wire [7:0] data_out22;
  output [7:0] data_out23;
  wire [7:0] data_out23;
  output [7:0] data_out24;
  wire [7:0] data_out24;
  output [7:0] data_out25;
  wire [7:0] data_out25;
  output [7:0] data_out26;
  wire [7:0] data_out26;
  output [7:0] data_out27;
  wire [7:0] data_out27;
  output [7:0] data_out28;
  wire [7:0] data_out28;
  output [7:0] data_out29;
  wire [7:0] data_out29;
  output [7:0] data_out30;
  wire [7:0] data_out30;
  output [7:0] data_out33;
  wire [7:0] data_out33;
  output [7:0] data_out34;
  wire [7:0] data_out34;
  output [7:0] data_out35;
  wire [7:0] data_out35;
  output [7:0] data_out36;
  wire [7:0] data_out36;
  output [7:0] data_out37;
  wire [7:0] data_out37;
  output [7:0] data_out38;
  wire [7:0] data_out38;
  output [7:0] data_out39;
  wire [7:0] data_out39;
  output [7:0] data_out40;
  wire [7:0] data_out40;
  output [7:0] data_out41;
  wire [7:0] data_out41;
  output [7:0] data_out42;
  wire [7:0] data_out42;
  output [7:0] data_out43;
  wire [7:0] data_out43;
  output [7:0] data_out44;
  wire [7:0] data_out44;
  output [7:0] data_out45;
  wire [7:0] data_out45;
  output [7:0] data_out46;
  wire [7:0] data_out46;
  output [7:0] data_out49;
  wire [7:0] data_out49;
  output [7:0] data_out50;
  wire [7:0] data_out50;
  output [7:0] data_out51;
  wire [7:0] data_out51;
  output [7:0] data_out52;
  wire [7:0] data_out52;
  output [7:0] data_out53;
  wire [7:0] data_out53;
  output [7:0] data_out54;
  wire [7:0] data_out54;
  output [7:0] data_out55;
  wire [7:0] data_out55;
  output [7:0] data_out56;
  wire [7:0] data_out56;
  output [7:0] data_out57;
  wire [7:0] data_out57;
  output [7:0] data_out58;
  wire [7:0] data_out58;
  output [7:0] data_out59;
  wire [7:0] data_out59;
  output [7:0] data_out60;
  wire [7:0] data_out60;
  output [7:0] data_out61;
  wire [7:0] data_out61;
  output [7:0] data_out62;
  wire [7:0] data_out62;
  output [7:0] data_out65;
  wire [7:0] data_out65;
  output [7:0] data_out66;
  wire [7:0] data_out66;
  output [7:0] data_out67;
  wire [7:0] data_out67;
  output [7:0] data_out68;
  wire [7:0] data_out68;
  output [7:0] data_out69;
  wire [7:0] data_out69;
  output [7:0] data_out70;
  wire [7:0] data_out70;
  output [7:0] data_out71;
  wire [7:0] data_out71;
  output [7:0] data_out72;
  wire [7:0] data_out72;
  output [7:0] data_out73;
  wire [7:0] data_out73;
  output [7:0] data_out74;
  wire [7:0] data_out74;
  output [7:0] data_out75;
  wire [7:0] data_out75;
  output [7:0] data_out76;
  wire [7:0] data_out76;
  output [7:0] data_out77;
  wire [7:0] data_out77;
  output [7:0] data_out78;
  wire [7:0] data_out78;
  output [7:0] data_out81;
  wire [7:0] data_out81;
  output [7:0] data_out82;
  wire [7:0] data_out82;
  output [7:0] data_out83;
  wire [7:0] data_out83;
  output [7:0] data_out84;
  wire [7:0] data_out84;
  output [7:0] data_out85;
  wire [7:0] data_out85;
  output [7:0] data_out86;
  wire [7:0] data_out86;
  output [7:0] data_out87;
  wire [7:0] data_out87;
  output [7:0] data_out88;
  wire [7:0] data_out88;
  output [7:0] data_out89;
  wire [7:0] data_out89;
  output [7:0] data_out90;
  wire [7:0] data_out90;
  output [7:0] data_out91;
  wire [7:0] data_out91;
  output [7:0] data_out92;
  wire [7:0] data_out92;
  output [7:0] data_out93;
  wire [7:0] data_out93;
  output [7:0] data_out94;
  wire [7:0] data_out94;
  output [7:0] data_out97;
  wire [7:0] data_out97;
  output [7:0] data_out98;
  wire [7:0] data_out98;
  output [7:0] data_out99;
  wire [7:0] data_out99;
  output [7:0] data_out100;
  wire [7:0] data_out100;
  output [7:0] data_out101;
  wire [7:0] data_out101;
  output [7:0] data_out102;
  wire [7:0] data_out102;
  output [7:0] data_out103;
  wire [7:0] data_out103;
  output [7:0] data_out104;
  wire [7:0] data_out104;
  output [7:0] data_out105;
  wire [7:0] data_out105;
  output [7:0] data_out106;
  wire [7:0] data_out106;
  output [7:0] data_out107;
  wire [7:0] data_out107;
  output [7:0] data_out108;
  wire [7:0] data_out108;
  output [7:0] data_out109;
  wire [7:0] data_out109;
  output [7:0] data_out110;
  wire [7:0] data_out110;
  output [7:0] data_out_index17;
  wire [7:0] data_out_index17;
  output [7:0] data_out_index18;
  wire [7:0] data_out_index18;
  output [7:0] data_out_index19;
  wire [7:0] data_out_index19;
  output [7:0] data_out_index20;
  wire [7:0] data_out_index20;
  output [7:0] data_out_index21;
  wire [7:0] data_out_index21;
  output [7:0] data_out_index22;
  wire [7:0] data_out_index22;
  output [7:0] data_out_index23;
  wire [7:0] data_out_index23;
  output [7:0] data_out_index24;
  wire [7:0] data_out_index24;
  output [7:0] data_out_index25;
  wire [7:0] data_out_index25;
  output [7:0] data_out_index26;
  wire [7:0] data_out_index26;
  output [7:0] data_out_index27;
  wire [7:0] data_out_index27;
  output [7:0] data_out_index28;
  wire [7:0] data_out_index28;
  output [7:0] data_out_index29;
  wire [7:0] data_out_index29;
  output [7:0] data_out_index30;
  wire [7:0] data_out_index30;
  output [7:0] data_out_index33;
  wire [7:0] data_out_index33;
  output [7:0] data_out_index34;
  wire [7:0] data_out_index34;
  output [7:0] data_out_index35;
  wire [7:0] data_out_index35;
  output [7:0] data_out_index36;
  wire [7:0] data_out_index36;
  output [7:0] data_out_index37;
  wire [7:0] data_out_index37;
  output [7:0] data_out_index38;
  wire [7:0] data_out_index38;
  output [7:0] data_out_index39;
  wire [7:0] data_out_index39;
  output [7:0] data_out_index40;
  wire [7:0] data_out_index40;
  output [7:0] data_out_index41;
  wire [7:0] data_out_index41;
  output [7:0] data_out_index42;
  wire [7:0] data_out_index42;
  output [7:0] data_out_index43;
  wire [7:0] data_out_index43;
  output [7:0] data_out_index44;
  wire [7:0] data_out_index44;
  output [7:0] data_out_index45;
  wire [7:0] data_out_index45;
  output [7:0] data_out_index46;
  wire [7:0] data_out_index46;
  output [7:0] data_out_index49;
  wire [7:0] data_out_index49;
  output [7:0] data_out_index50;
  wire [7:0] data_out_index50;
  output [7:0] data_out_index51;
  wire [7:0] data_out_index51;
  output [7:0] data_out_index52;
  wire [7:0] data_out_index52;
  output [7:0] data_out_index53;
  wire [7:0] data_out_index53;
  output [7:0] data_out_index54;
  wire [7:0] data_out_index54;
  output [7:0] data_out_index55;
  wire [7:0] data_out_index55;
  output [7:0] data_out_index56;
  wire [7:0] data_out_index56;
  output [7:0] data_out_index57;
  wire [7:0] data_out_index57;
  output [7:0] data_out_index58;
  wire [7:0] data_out_index58;
  output [7:0] data_out_index59;
  wire [7:0] data_out_index59;
  output [7:0] data_out_index60;
  wire [7:0] data_out_index60;
  output [7:0] data_out_index61;
  wire [7:0] data_out_index61;
  output [7:0] data_out_index62;
  wire [7:0] data_out_index62;
  output [7:0] data_out_index65;
  wire [7:0] data_out_index65;
  output [7:0] data_out_index66;
  wire [7:0] data_out_index66;
  output [7:0] data_out_index67;
  wire [7:0] data_out_index67;
  output [7:0] data_out_index68;
  wire [7:0] data_out_index68;
  output [7:0] data_out_index69;
  wire [7:0] data_out_index69;
  output [7:0] data_out_index70;
  wire [7:0] data_out_index70;
  output [7:0] data_out_index71;
  wire [7:0] data_out_index71;
  output [7:0] data_out_index72;
  wire [7:0] data_out_index72;
  output [7:0] data_out_index73;
  wire [7:0] data_out_index73;
  output [7:0] data_out_index74;
  wire [7:0] data_out_index74;
  output [7:0] data_out_index75;
  wire [7:0] data_out_index75;
  output [7:0] data_out_index76;
  wire [7:0] data_out_index76;
  output [7:0] data_out_index77;
  wire [7:0] data_out_index77;
  output [7:0] data_out_index78;
  wire [7:0] data_out_index78;
  output [7:0] data_out_index81;
  wire [7:0] data_out_index81;
  output [7:0] data_out_index82;
  wire [7:0] data_out_index82;
  output [7:0] data_out_index83;
  wire [7:0] data_out_index83;
  output [7:0] data_out_index84;
  wire [7:0] data_out_index84;
  output [7:0] data_out_index85;
  wire [7:0] data_out_index85;
  output [7:0] data_out_index86;
  wire [7:0] data_out_index86;
  output [7:0] data_out_index87;
  wire [7:0] data_out_index87;
  output [7:0] data_out_index88;
  wire [7:0] data_out_index88;
  output [7:0] data_out_index89;
  wire [7:0] data_out_index89;
  output [7:0] data_out_index90;
  wire [7:0] data_out_index90;
  output [7:0] data_out_index91;
  wire [7:0] data_out_index91;
  output [7:0] data_out_index92;
  wire [7:0] data_out_index92;
  output [7:0] data_out_index93;
  wire [7:0] data_out_index93;
  output [7:0] data_out_index94;
  wire [7:0] data_out_index94;
  output [7:0] data_out_index97;
  wire [7:0] data_out_index97;
  output [7:0] data_out_index98;
  wire [7:0] data_out_index98;
  output [7:0] data_out_index99;
  wire [7:0] data_out_index99;
  output [7:0] data_out_index100;
  wire [7:0] data_out_index100;
  output [7:0] data_out_index101;
  wire [7:0] data_out_index101;
  output [7:0] data_out_index102;
  wire [7:0] data_out_index102;
  output [7:0] data_out_index103;
  wire [7:0] data_out_index103;
  output [7:0] data_out_index104;
  wire [7:0] data_out_index104;
  output [7:0] data_out_index105;
  wire [7:0] data_out_index105;
  output [7:0] data_out_index106;
  wire [7:0] data_out_index106;
  output [7:0] data_out_index107;
  wire [7:0] data_out_index107;
  output [7:0] data_out_index108;
  wire [7:0] data_out_index108;
  output [7:0] data_out_index109;
  wire [7:0] data_out_index109;
  output [7:0] data_out_index110;
  wire [7:0] data_out_index110;
  input [7:0] distance_count_all;
  wire [7:0] distance_count_all;
  output [127:0] all_sg_out17;
  wire [127:0] all_sg_out17;
  output [127:0] all_sg_out18;
  wire [127:0] all_sg_out18;
  output [127:0] all_sg_out19;
  wire [127:0] all_sg_out19;
  output [127:0] all_sg_out20;
  wire [127:0] all_sg_out20;
  output [127:0] all_sg_out21;
  wire [127:0] all_sg_out21;
  output [127:0] all_sg_out22;
  wire [127:0] all_sg_out22;
  output [127:0] all_sg_out23;
  wire [127:0] all_sg_out23;
  output [127:0] all_sg_out24;
  wire [127:0] all_sg_out24;
  output [127:0] all_sg_out25;
  wire [127:0] all_sg_out25;
  output [127:0] all_sg_out26;
  wire [127:0] all_sg_out26;
  output [127:0] all_sg_out27;
  wire [127:0] all_sg_out27;
  output [127:0] all_sg_out28;
  wire [127:0] all_sg_out28;
  output [127:0] all_sg_out29;
  wire [127:0] all_sg_out29;
  output [127:0] all_sg_out30;
  wire [127:0] all_sg_out30;
  output [127:0] all_sg_out33;
  wire [127:0] all_sg_out33;
  output [127:0] all_sg_out34;
  wire [127:0] all_sg_out34;
  output [127:0] all_sg_out35;
  wire [127:0] all_sg_out35;
  output [127:0] all_sg_out36;
  wire [127:0] all_sg_out36;
  output [127:0] all_sg_out37;
  wire [127:0] all_sg_out37;
  output [127:0] all_sg_out38;
  wire [127:0] all_sg_out38;
  output [127:0] all_sg_out39;
  wire [127:0] all_sg_out39;
  output [127:0] all_sg_out40;
  wire [127:0] all_sg_out40;
  output [127:0] all_sg_out41;
  wire [127:0] all_sg_out41;
  output [127:0] all_sg_out42;
  wire [127:0] all_sg_out42;
  output [127:0] all_sg_out43;
  wire [127:0] all_sg_out43;
  output [127:0] all_sg_out44;
  wire [127:0] all_sg_out44;
  output [127:0] all_sg_out45;
  wire [127:0] all_sg_out45;
  output [127:0] all_sg_out46;
  wire [127:0] all_sg_out46;
  output [127:0] all_sg_out49;
  wire [127:0] all_sg_out49;
  output [127:0] all_sg_out50;
  wire [127:0] all_sg_out50;
  output [127:0] all_sg_out51;
  wire [127:0] all_sg_out51;
  output [127:0] all_sg_out52;
  wire [127:0] all_sg_out52;
  output [127:0] all_sg_out53;
  wire [127:0] all_sg_out53;
  output [127:0] all_sg_out54;
  wire [127:0] all_sg_out54;
  output [127:0] all_sg_out55;
  wire [127:0] all_sg_out55;
  output [127:0] all_sg_out56;
  wire [127:0] all_sg_out56;
  output [127:0] all_sg_out57;
  wire [127:0] all_sg_out57;
  output [127:0] all_sg_out58;
  wire [127:0] all_sg_out58;
  output [127:0] all_sg_out59;
  wire [127:0] all_sg_out59;
  output [127:0] all_sg_out60;
  wire [127:0] all_sg_out60;
  output [127:0] all_sg_out61;
  wire [127:0] all_sg_out61;
  output [127:0] all_sg_out62;
  wire [127:0] all_sg_out62;
  output [127:0] all_sg_out65;
  wire [127:0] all_sg_out65;
  output [127:0] all_sg_out66;
  wire [127:0] all_sg_out66;
  output [127:0] all_sg_out67;
  wire [127:0] all_sg_out67;
  output [127:0] all_sg_out68;
  wire [127:0] all_sg_out68;
  output [127:0] all_sg_out69;
  wire [127:0] all_sg_out69;
  output [127:0] all_sg_out70;
  wire [127:0] all_sg_out70;
  output [127:0] all_sg_out71;
  wire [127:0] all_sg_out71;
  output [127:0] all_sg_out72;
  wire [127:0] all_sg_out72;
  output [127:0] all_sg_out73;
  wire [127:0] all_sg_out73;
  output [127:0] all_sg_out74;
  wire [127:0] all_sg_out74;
  output [127:0] all_sg_out75;
  wire [127:0] all_sg_out75;
  output [127:0] all_sg_out76;
  wire [127:0] all_sg_out76;
  output [127:0] all_sg_out77;
  wire [127:0] all_sg_out77;
  output [127:0] all_sg_out78;
  wire [127:0] all_sg_out78;
  output [127:0] all_sg_out81;
  wire [127:0] all_sg_out81;
  output [127:0] all_sg_out82;
  wire [127:0] all_sg_out82;
  output [127:0] all_sg_out83;
  wire [127:0] all_sg_out83;
  output [127:0] all_sg_out84;
  wire [127:0] all_sg_out84;
  output [127:0] all_sg_out85;
  wire [127:0] all_sg_out85;
  output [127:0] all_sg_out86;
  wire [127:0] all_sg_out86;
  output [127:0] all_sg_out87;
  wire [127:0] all_sg_out87;
  output [127:0] all_sg_out88;
  wire [127:0] all_sg_out88;
  output [127:0] all_sg_out89;
  wire [127:0] all_sg_out89;
  output [127:0] all_sg_out90;
  wire [127:0] all_sg_out90;
  output [127:0] all_sg_out91;
  wire [127:0] all_sg_out91;
  output [127:0] all_sg_out92;
  wire [127:0] all_sg_out92;
  output [127:0] all_sg_out93;
  wire [127:0] all_sg_out93;
  output [127:0] all_sg_out94;
  wire [127:0] all_sg_out94;
  output [127:0] all_sg_out97;
  wire [127:0] all_sg_out97;
  output [127:0] all_sg_out98;
  wire [127:0] all_sg_out98;
  output [127:0] all_sg_out99;
  wire [127:0] all_sg_out99;
  output [127:0] all_sg_out100;
  wire [127:0] all_sg_out100;
  output [127:0] all_sg_out101;
  wire [127:0] all_sg_out101;
  output [127:0] all_sg_out102;
  wire [127:0] all_sg_out102;
  output [127:0] all_sg_out103;
  wire [127:0] all_sg_out103;
  output [127:0] all_sg_out104;
  wire [127:0] all_sg_out104;
  output [127:0] all_sg_out105;
  wire [127:0] all_sg_out105;
  output [127:0] all_sg_out106;
  wire [127:0] all_sg_out106;
  output [127:0] all_sg_out107;
  wire [127:0] all_sg_out107;
  output [127:0] all_sg_out108;
  wire [127:0] all_sg_out108;
  output [127:0] all_sg_out109;
  wire [127:0] all_sg_out109;
  output [127:0] all_sg_out110;
  wire [127:0] all_sg_out110;
  input in_do;
  wire in_do;
  output out_do;
  wire out_do;
  output out_data;
  wire out_data;
  wire dig_add_all;
  reg sig_reg;
  wire [127:0] _add_map_x_wall_end_in;
  wire [127:0] _add_map_x_all_sg_up;
  wire [127:0] _add_map_x_all_sg_down;
  wire [127:0] _add_map_x_all_sg_right;
  wire [127:0] _add_map_x_all_sg_left;
  wire [7:0] _add_map_x_moto_org_near;
  wire [7:0] _add_map_x_moto_org_near1;
  wire [7:0] _add_map_x_moto_org_near2;
  wire [7:0] _add_map_x_moto_org_near3;
  wire [7:0] _add_map_x_moto_org;
  wire [1:0] _add_map_x_sg_up;
  wire [1:0] _add_map_x_sg_down;
  wire [1:0] _add_map_x_sg_left;
  wire [1:0] _add_map_x_sg_right;
  wire _add_map_x_wall_t_in;
  wire [7:0] _add_map_x_moto;
  wire [7:0] _add_map_x_up;
  wire [7:0] _add_map_x_right;
  wire [7:0] _add_map_x_down;
  wire [7:0] _add_map_x_left;
  wire [7:0] _add_map_x_start;
  wire [7:0] _add_map_x_goal;
  wire [7:0] _add_map_x_now;
  wire [7:0] _add_map_x_distance;
  wire [127:0] _add_map_x_end_wall;
  wire [127:0] _add_map_x_all_s_g;
  wire [127:0] _add_map_x_all_s_g_near;
  wire [7:0] _add_map_x_data_out;
  wire [7:0] _add_map_x_data_out_index;
  wire [7:0] _add_map_x_data_near;
  wire _add_map_x_wall_t_out;
  wire [7:0] _add_map_x_data_org;
  wire [7:0] _add_map_x_data_org_near;
  wire [1:0] _add_map_x_s_g;
  wire [1:0] _add_map_x_s_g_near;
  wire _add_map_x_add_exe;
  wire _add_map_x_p_reset;
  wire _add_map_x_m_clock;
  wire [127:0] _add_map_x_41_wall_end_in;
  wire [127:0] _add_map_x_41_all_sg_up;
  wire [127:0] _add_map_x_41_all_sg_down;
  wire [127:0] _add_map_x_41_all_sg_right;
  wire [127:0] _add_map_x_41_all_sg_left;
  wire [7:0] _add_map_x_41_moto_org_near;
  wire [7:0] _add_map_x_41_moto_org_near1;
  wire [7:0] _add_map_x_41_moto_org_near2;
  wire [7:0] _add_map_x_41_moto_org_near3;
  wire [7:0] _add_map_x_41_moto_org;
  wire [1:0] _add_map_x_41_sg_up;
  wire [1:0] _add_map_x_41_sg_down;
  wire [1:0] _add_map_x_41_sg_left;
  wire [1:0] _add_map_x_41_sg_right;
  wire _add_map_x_41_wall_t_in;
  wire [7:0] _add_map_x_41_moto;
  wire [7:0] _add_map_x_41_up;
  wire [7:0] _add_map_x_41_right;
  wire [7:0] _add_map_x_41_down;
  wire [7:0] _add_map_x_41_left;
  wire [7:0] _add_map_x_41_start;
  wire [7:0] _add_map_x_41_goal;
  wire [7:0] _add_map_x_41_now;
  wire [7:0] _add_map_x_41_distance;
  wire [127:0] _add_map_x_41_end_wall;
  wire [127:0] _add_map_x_41_all_s_g;
  wire [127:0] _add_map_x_41_all_s_g_near;
  wire [7:0] _add_map_x_41_data_out;
  wire [7:0] _add_map_x_41_data_out_index;
  wire [7:0] _add_map_x_41_data_near;
  wire _add_map_x_41_wall_t_out;
  wire [7:0] _add_map_x_41_data_org;
  wire [7:0] _add_map_x_41_data_org_near;
  wire [1:0] _add_map_x_41_s_g;
  wire [1:0] _add_map_x_41_s_g_near;
  wire _add_map_x_41_add_exe;
  wire _add_map_x_41_p_reset;
  wire _add_map_x_41_m_clock;
  wire [127:0] _add_map_x_40_wall_end_in;
  wire [127:0] _add_map_x_40_all_sg_up;
  wire [127:0] _add_map_x_40_all_sg_down;
  wire [127:0] _add_map_x_40_all_sg_right;
  wire [127:0] _add_map_x_40_all_sg_left;
  wire [7:0] _add_map_x_40_moto_org_near;
  wire [7:0] _add_map_x_40_moto_org_near1;
  wire [7:0] _add_map_x_40_moto_org_near2;
  wire [7:0] _add_map_x_40_moto_org_near3;
  wire [7:0] _add_map_x_40_moto_org;
  wire [1:0] _add_map_x_40_sg_up;
  wire [1:0] _add_map_x_40_sg_down;
  wire [1:0] _add_map_x_40_sg_left;
  wire [1:0] _add_map_x_40_sg_right;
  wire _add_map_x_40_wall_t_in;
  wire [7:0] _add_map_x_40_moto;
  wire [7:0] _add_map_x_40_up;
  wire [7:0] _add_map_x_40_right;
  wire [7:0] _add_map_x_40_down;
  wire [7:0] _add_map_x_40_left;
  wire [7:0] _add_map_x_40_start;
  wire [7:0] _add_map_x_40_goal;
  wire [7:0] _add_map_x_40_now;
  wire [7:0] _add_map_x_40_distance;
  wire [127:0] _add_map_x_40_end_wall;
  wire [127:0] _add_map_x_40_all_s_g;
  wire [127:0] _add_map_x_40_all_s_g_near;
  wire [7:0] _add_map_x_40_data_out;
  wire [7:0] _add_map_x_40_data_out_index;
  wire [7:0] _add_map_x_40_data_near;
  wire _add_map_x_40_wall_t_out;
  wire [7:0] _add_map_x_40_data_org;
  wire [7:0] _add_map_x_40_data_org_near;
  wire [1:0] _add_map_x_40_s_g;
  wire [1:0] _add_map_x_40_s_g_near;
  wire _add_map_x_40_add_exe;
  wire _add_map_x_40_p_reset;
  wire _add_map_x_40_m_clock;
  wire [127:0] _add_map_x_39_wall_end_in;
  wire [127:0] _add_map_x_39_all_sg_up;
  wire [127:0] _add_map_x_39_all_sg_down;
  wire [127:0] _add_map_x_39_all_sg_right;
  wire [127:0] _add_map_x_39_all_sg_left;
  wire [7:0] _add_map_x_39_moto_org_near;
  wire [7:0] _add_map_x_39_moto_org_near1;
  wire [7:0] _add_map_x_39_moto_org_near2;
  wire [7:0] _add_map_x_39_moto_org_near3;
  wire [7:0] _add_map_x_39_moto_org;
  wire [1:0] _add_map_x_39_sg_up;
  wire [1:0] _add_map_x_39_sg_down;
  wire [1:0] _add_map_x_39_sg_left;
  wire [1:0] _add_map_x_39_sg_right;
  wire _add_map_x_39_wall_t_in;
  wire [7:0] _add_map_x_39_moto;
  wire [7:0] _add_map_x_39_up;
  wire [7:0] _add_map_x_39_right;
  wire [7:0] _add_map_x_39_down;
  wire [7:0] _add_map_x_39_left;
  wire [7:0] _add_map_x_39_start;
  wire [7:0] _add_map_x_39_goal;
  wire [7:0] _add_map_x_39_now;
  wire [7:0] _add_map_x_39_distance;
  wire [127:0] _add_map_x_39_end_wall;
  wire [127:0] _add_map_x_39_all_s_g;
  wire [127:0] _add_map_x_39_all_s_g_near;
  wire [7:0] _add_map_x_39_data_out;
  wire [7:0] _add_map_x_39_data_out_index;
  wire [7:0] _add_map_x_39_data_near;
  wire _add_map_x_39_wall_t_out;
  wire [7:0] _add_map_x_39_data_org;
  wire [7:0] _add_map_x_39_data_org_near;
  wire [1:0] _add_map_x_39_s_g;
  wire [1:0] _add_map_x_39_s_g_near;
  wire _add_map_x_39_add_exe;
  wire _add_map_x_39_p_reset;
  wire _add_map_x_39_m_clock;
  wire [127:0] _add_map_x_38_wall_end_in;
  wire [127:0] _add_map_x_38_all_sg_up;
  wire [127:0] _add_map_x_38_all_sg_down;
  wire [127:0] _add_map_x_38_all_sg_right;
  wire [127:0] _add_map_x_38_all_sg_left;
  wire [7:0] _add_map_x_38_moto_org_near;
  wire [7:0] _add_map_x_38_moto_org_near1;
  wire [7:0] _add_map_x_38_moto_org_near2;
  wire [7:0] _add_map_x_38_moto_org_near3;
  wire [7:0] _add_map_x_38_moto_org;
  wire [1:0] _add_map_x_38_sg_up;
  wire [1:0] _add_map_x_38_sg_down;
  wire [1:0] _add_map_x_38_sg_left;
  wire [1:0] _add_map_x_38_sg_right;
  wire _add_map_x_38_wall_t_in;
  wire [7:0] _add_map_x_38_moto;
  wire [7:0] _add_map_x_38_up;
  wire [7:0] _add_map_x_38_right;
  wire [7:0] _add_map_x_38_down;
  wire [7:0] _add_map_x_38_left;
  wire [7:0] _add_map_x_38_start;
  wire [7:0] _add_map_x_38_goal;
  wire [7:0] _add_map_x_38_now;
  wire [7:0] _add_map_x_38_distance;
  wire [127:0] _add_map_x_38_end_wall;
  wire [127:0] _add_map_x_38_all_s_g;
  wire [127:0] _add_map_x_38_all_s_g_near;
  wire [7:0] _add_map_x_38_data_out;
  wire [7:0] _add_map_x_38_data_out_index;
  wire [7:0] _add_map_x_38_data_near;
  wire _add_map_x_38_wall_t_out;
  wire [7:0] _add_map_x_38_data_org;
  wire [7:0] _add_map_x_38_data_org_near;
  wire [1:0] _add_map_x_38_s_g;
  wire [1:0] _add_map_x_38_s_g_near;
  wire _add_map_x_38_add_exe;
  wire _add_map_x_38_p_reset;
  wire _add_map_x_38_m_clock;
  wire [127:0] _add_map_x_37_wall_end_in;
  wire [127:0] _add_map_x_37_all_sg_up;
  wire [127:0] _add_map_x_37_all_sg_down;
  wire [127:0] _add_map_x_37_all_sg_right;
  wire [127:0] _add_map_x_37_all_sg_left;
  wire [7:0] _add_map_x_37_moto_org_near;
  wire [7:0] _add_map_x_37_moto_org_near1;
  wire [7:0] _add_map_x_37_moto_org_near2;
  wire [7:0] _add_map_x_37_moto_org_near3;
  wire [7:0] _add_map_x_37_moto_org;
  wire [1:0] _add_map_x_37_sg_up;
  wire [1:0] _add_map_x_37_sg_down;
  wire [1:0] _add_map_x_37_sg_left;
  wire [1:0] _add_map_x_37_sg_right;
  wire _add_map_x_37_wall_t_in;
  wire [7:0] _add_map_x_37_moto;
  wire [7:0] _add_map_x_37_up;
  wire [7:0] _add_map_x_37_right;
  wire [7:0] _add_map_x_37_down;
  wire [7:0] _add_map_x_37_left;
  wire [7:0] _add_map_x_37_start;
  wire [7:0] _add_map_x_37_goal;
  wire [7:0] _add_map_x_37_now;
  wire [7:0] _add_map_x_37_distance;
  wire [127:0] _add_map_x_37_end_wall;
  wire [127:0] _add_map_x_37_all_s_g;
  wire [127:0] _add_map_x_37_all_s_g_near;
  wire [7:0] _add_map_x_37_data_out;
  wire [7:0] _add_map_x_37_data_out_index;
  wire [7:0] _add_map_x_37_data_near;
  wire _add_map_x_37_wall_t_out;
  wire [7:0] _add_map_x_37_data_org;
  wire [7:0] _add_map_x_37_data_org_near;
  wire [1:0] _add_map_x_37_s_g;
  wire [1:0] _add_map_x_37_s_g_near;
  wire _add_map_x_37_add_exe;
  wire _add_map_x_37_p_reset;
  wire _add_map_x_37_m_clock;
  wire [127:0] _add_map_x_36_wall_end_in;
  wire [127:0] _add_map_x_36_all_sg_up;
  wire [127:0] _add_map_x_36_all_sg_down;
  wire [127:0] _add_map_x_36_all_sg_right;
  wire [127:0] _add_map_x_36_all_sg_left;
  wire [7:0] _add_map_x_36_moto_org_near;
  wire [7:0] _add_map_x_36_moto_org_near1;
  wire [7:0] _add_map_x_36_moto_org_near2;
  wire [7:0] _add_map_x_36_moto_org_near3;
  wire [7:0] _add_map_x_36_moto_org;
  wire [1:0] _add_map_x_36_sg_up;
  wire [1:0] _add_map_x_36_sg_down;
  wire [1:0] _add_map_x_36_sg_left;
  wire [1:0] _add_map_x_36_sg_right;
  wire _add_map_x_36_wall_t_in;
  wire [7:0] _add_map_x_36_moto;
  wire [7:0] _add_map_x_36_up;
  wire [7:0] _add_map_x_36_right;
  wire [7:0] _add_map_x_36_down;
  wire [7:0] _add_map_x_36_left;
  wire [7:0] _add_map_x_36_start;
  wire [7:0] _add_map_x_36_goal;
  wire [7:0] _add_map_x_36_now;
  wire [7:0] _add_map_x_36_distance;
  wire [127:0] _add_map_x_36_end_wall;
  wire [127:0] _add_map_x_36_all_s_g;
  wire [127:0] _add_map_x_36_all_s_g_near;
  wire [7:0] _add_map_x_36_data_out;
  wire [7:0] _add_map_x_36_data_out_index;
  wire [7:0] _add_map_x_36_data_near;
  wire _add_map_x_36_wall_t_out;
  wire [7:0] _add_map_x_36_data_org;
  wire [7:0] _add_map_x_36_data_org_near;
  wire [1:0] _add_map_x_36_s_g;
  wire [1:0] _add_map_x_36_s_g_near;
  wire _add_map_x_36_add_exe;
  wire _add_map_x_36_p_reset;
  wire _add_map_x_36_m_clock;
  wire [127:0] _add_map_x_35_wall_end_in;
  wire [127:0] _add_map_x_35_all_sg_up;
  wire [127:0] _add_map_x_35_all_sg_down;
  wire [127:0] _add_map_x_35_all_sg_right;
  wire [127:0] _add_map_x_35_all_sg_left;
  wire [7:0] _add_map_x_35_moto_org_near;
  wire [7:0] _add_map_x_35_moto_org_near1;
  wire [7:0] _add_map_x_35_moto_org_near2;
  wire [7:0] _add_map_x_35_moto_org_near3;
  wire [7:0] _add_map_x_35_moto_org;
  wire [1:0] _add_map_x_35_sg_up;
  wire [1:0] _add_map_x_35_sg_down;
  wire [1:0] _add_map_x_35_sg_left;
  wire [1:0] _add_map_x_35_sg_right;
  wire _add_map_x_35_wall_t_in;
  wire [7:0] _add_map_x_35_moto;
  wire [7:0] _add_map_x_35_up;
  wire [7:0] _add_map_x_35_right;
  wire [7:0] _add_map_x_35_down;
  wire [7:0] _add_map_x_35_left;
  wire [7:0] _add_map_x_35_start;
  wire [7:0] _add_map_x_35_goal;
  wire [7:0] _add_map_x_35_now;
  wire [7:0] _add_map_x_35_distance;
  wire [127:0] _add_map_x_35_end_wall;
  wire [127:0] _add_map_x_35_all_s_g;
  wire [127:0] _add_map_x_35_all_s_g_near;
  wire [7:0] _add_map_x_35_data_out;
  wire [7:0] _add_map_x_35_data_out_index;
  wire [7:0] _add_map_x_35_data_near;
  wire _add_map_x_35_wall_t_out;
  wire [7:0] _add_map_x_35_data_org;
  wire [7:0] _add_map_x_35_data_org_near;
  wire [1:0] _add_map_x_35_s_g;
  wire [1:0] _add_map_x_35_s_g_near;
  wire _add_map_x_35_add_exe;
  wire _add_map_x_35_p_reset;
  wire _add_map_x_35_m_clock;
  wire [127:0] _add_map_x_34_wall_end_in;
  wire [127:0] _add_map_x_34_all_sg_up;
  wire [127:0] _add_map_x_34_all_sg_down;
  wire [127:0] _add_map_x_34_all_sg_right;
  wire [127:0] _add_map_x_34_all_sg_left;
  wire [7:0] _add_map_x_34_moto_org_near;
  wire [7:0] _add_map_x_34_moto_org_near1;
  wire [7:0] _add_map_x_34_moto_org_near2;
  wire [7:0] _add_map_x_34_moto_org_near3;
  wire [7:0] _add_map_x_34_moto_org;
  wire [1:0] _add_map_x_34_sg_up;
  wire [1:0] _add_map_x_34_sg_down;
  wire [1:0] _add_map_x_34_sg_left;
  wire [1:0] _add_map_x_34_sg_right;
  wire _add_map_x_34_wall_t_in;
  wire [7:0] _add_map_x_34_moto;
  wire [7:0] _add_map_x_34_up;
  wire [7:0] _add_map_x_34_right;
  wire [7:0] _add_map_x_34_down;
  wire [7:0] _add_map_x_34_left;
  wire [7:0] _add_map_x_34_start;
  wire [7:0] _add_map_x_34_goal;
  wire [7:0] _add_map_x_34_now;
  wire [7:0] _add_map_x_34_distance;
  wire [127:0] _add_map_x_34_end_wall;
  wire [127:0] _add_map_x_34_all_s_g;
  wire [127:0] _add_map_x_34_all_s_g_near;
  wire [7:0] _add_map_x_34_data_out;
  wire [7:0] _add_map_x_34_data_out_index;
  wire [7:0] _add_map_x_34_data_near;
  wire _add_map_x_34_wall_t_out;
  wire [7:0] _add_map_x_34_data_org;
  wire [7:0] _add_map_x_34_data_org_near;
  wire [1:0] _add_map_x_34_s_g;
  wire [1:0] _add_map_x_34_s_g_near;
  wire _add_map_x_34_add_exe;
  wire _add_map_x_34_p_reset;
  wire _add_map_x_34_m_clock;
  wire [127:0] _add_map_x_33_wall_end_in;
  wire [127:0] _add_map_x_33_all_sg_up;
  wire [127:0] _add_map_x_33_all_sg_down;
  wire [127:0] _add_map_x_33_all_sg_right;
  wire [127:0] _add_map_x_33_all_sg_left;
  wire [7:0] _add_map_x_33_moto_org_near;
  wire [7:0] _add_map_x_33_moto_org_near1;
  wire [7:0] _add_map_x_33_moto_org_near2;
  wire [7:0] _add_map_x_33_moto_org_near3;
  wire [7:0] _add_map_x_33_moto_org;
  wire [1:0] _add_map_x_33_sg_up;
  wire [1:0] _add_map_x_33_sg_down;
  wire [1:0] _add_map_x_33_sg_left;
  wire [1:0] _add_map_x_33_sg_right;
  wire _add_map_x_33_wall_t_in;
  wire [7:0] _add_map_x_33_moto;
  wire [7:0] _add_map_x_33_up;
  wire [7:0] _add_map_x_33_right;
  wire [7:0] _add_map_x_33_down;
  wire [7:0] _add_map_x_33_left;
  wire [7:0] _add_map_x_33_start;
  wire [7:0] _add_map_x_33_goal;
  wire [7:0] _add_map_x_33_now;
  wire [7:0] _add_map_x_33_distance;
  wire [127:0] _add_map_x_33_end_wall;
  wire [127:0] _add_map_x_33_all_s_g;
  wire [127:0] _add_map_x_33_all_s_g_near;
  wire [7:0] _add_map_x_33_data_out;
  wire [7:0] _add_map_x_33_data_out_index;
  wire [7:0] _add_map_x_33_data_near;
  wire _add_map_x_33_wall_t_out;
  wire [7:0] _add_map_x_33_data_org;
  wire [7:0] _add_map_x_33_data_org_near;
  wire [1:0] _add_map_x_33_s_g;
  wire [1:0] _add_map_x_33_s_g_near;
  wire _add_map_x_33_add_exe;
  wire _add_map_x_33_p_reset;
  wire _add_map_x_33_m_clock;
  wire [127:0] _add_map_x_32_wall_end_in;
  wire [127:0] _add_map_x_32_all_sg_up;
  wire [127:0] _add_map_x_32_all_sg_down;
  wire [127:0] _add_map_x_32_all_sg_right;
  wire [127:0] _add_map_x_32_all_sg_left;
  wire [7:0] _add_map_x_32_moto_org_near;
  wire [7:0] _add_map_x_32_moto_org_near1;
  wire [7:0] _add_map_x_32_moto_org_near2;
  wire [7:0] _add_map_x_32_moto_org_near3;
  wire [7:0] _add_map_x_32_moto_org;
  wire [1:0] _add_map_x_32_sg_up;
  wire [1:0] _add_map_x_32_sg_down;
  wire [1:0] _add_map_x_32_sg_left;
  wire [1:0] _add_map_x_32_sg_right;
  wire _add_map_x_32_wall_t_in;
  wire [7:0] _add_map_x_32_moto;
  wire [7:0] _add_map_x_32_up;
  wire [7:0] _add_map_x_32_right;
  wire [7:0] _add_map_x_32_down;
  wire [7:0] _add_map_x_32_left;
  wire [7:0] _add_map_x_32_start;
  wire [7:0] _add_map_x_32_goal;
  wire [7:0] _add_map_x_32_now;
  wire [7:0] _add_map_x_32_distance;
  wire [127:0] _add_map_x_32_end_wall;
  wire [127:0] _add_map_x_32_all_s_g;
  wire [127:0] _add_map_x_32_all_s_g_near;
  wire [7:0] _add_map_x_32_data_out;
  wire [7:0] _add_map_x_32_data_out_index;
  wire [7:0] _add_map_x_32_data_near;
  wire _add_map_x_32_wall_t_out;
  wire [7:0] _add_map_x_32_data_org;
  wire [7:0] _add_map_x_32_data_org_near;
  wire [1:0] _add_map_x_32_s_g;
  wire [1:0] _add_map_x_32_s_g_near;
  wire _add_map_x_32_add_exe;
  wire _add_map_x_32_p_reset;
  wire _add_map_x_32_m_clock;
  wire [127:0] _add_map_x_31_wall_end_in;
  wire [127:0] _add_map_x_31_all_sg_up;
  wire [127:0] _add_map_x_31_all_sg_down;
  wire [127:0] _add_map_x_31_all_sg_right;
  wire [127:0] _add_map_x_31_all_sg_left;
  wire [7:0] _add_map_x_31_moto_org_near;
  wire [7:0] _add_map_x_31_moto_org_near1;
  wire [7:0] _add_map_x_31_moto_org_near2;
  wire [7:0] _add_map_x_31_moto_org_near3;
  wire [7:0] _add_map_x_31_moto_org;
  wire [1:0] _add_map_x_31_sg_up;
  wire [1:0] _add_map_x_31_sg_down;
  wire [1:0] _add_map_x_31_sg_left;
  wire [1:0] _add_map_x_31_sg_right;
  wire _add_map_x_31_wall_t_in;
  wire [7:0] _add_map_x_31_moto;
  wire [7:0] _add_map_x_31_up;
  wire [7:0] _add_map_x_31_right;
  wire [7:0] _add_map_x_31_down;
  wire [7:0] _add_map_x_31_left;
  wire [7:0] _add_map_x_31_start;
  wire [7:0] _add_map_x_31_goal;
  wire [7:0] _add_map_x_31_now;
  wire [7:0] _add_map_x_31_distance;
  wire [127:0] _add_map_x_31_end_wall;
  wire [127:0] _add_map_x_31_all_s_g;
  wire [127:0] _add_map_x_31_all_s_g_near;
  wire [7:0] _add_map_x_31_data_out;
  wire [7:0] _add_map_x_31_data_out_index;
  wire [7:0] _add_map_x_31_data_near;
  wire _add_map_x_31_wall_t_out;
  wire [7:0] _add_map_x_31_data_org;
  wire [7:0] _add_map_x_31_data_org_near;
  wire [1:0] _add_map_x_31_s_g;
  wire [1:0] _add_map_x_31_s_g_near;
  wire _add_map_x_31_add_exe;
  wire _add_map_x_31_p_reset;
  wire _add_map_x_31_m_clock;
  wire [127:0] _add_map_x_30_wall_end_in;
  wire [127:0] _add_map_x_30_all_sg_up;
  wire [127:0] _add_map_x_30_all_sg_down;
  wire [127:0] _add_map_x_30_all_sg_right;
  wire [127:0] _add_map_x_30_all_sg_left;
  wire [7:0] _add_map_x_30_moto_org_near;
  wire [7:0] _add_map_x_30_moto_org_near1;
  wire [7:0] _add_map_x_30_moto_org_near2;
  wire [7:0] _add_map_x_30_moto_org_near3;
  wire [7:0] _add_map_x_30_moto_org;
  wire [1:0] _add_map_x_30_sg_up;
  wire [1:0] _add_map_x_30_sg_down;
  wire [1:0] _add_map_x_30_sg_left;
  wire [1:0] _add_map_x_30_sg_right;
  wire _add_map_x_30_wall_t_in;
  wire [7:0] _add_map_x_30_moto;
  wire [7:0] _add_map_x_30_up;
  wire [7:0] _add_map_x_30_right;
  wire [7:0] _add_map_x_30_down;
  wire [7:0] _add_map_x_30_left;
  wire [7:0] _add_map_x_30_start;
  wire [7:0] _add_map_x_30_goal;
  wire [7:0] _add_map_x_30_now;
  wire [7:0] _add_map_x_30_distance;
  wire [127:0] _add_map_x_30_end_wall;
  wire [127:0] _add_map_x_30_all_s_g;
  wire [127:0] _add_map_x_30_all_s_g_near;
  wire [7:0] _add_map_x_30_data_out;
  wire [7:0] _add_map_x_30_data_out_index;
  wire [7:0] _add_map_x_30_data_near;
  wire _add_map_x_30_wall_t_out;
  wire [7:0] _add_map_x_30_data_org;
  wire [7:0] _add_map_x_30_data_org_near;
  wire [1:0] _add_map_x_30_s_g;
  wire [1:0] _add_map_x_30_s_g_near;
  wire _add_map_x_30_add_exe;
  wire _add_map_x_30_p_reset;
  wire _add_map_x_30_m_clock;
  wire [127:0] _add_map_x_29_wall_end_in;
  wire [127:0] _add_map_x_29_all_sg_up;
  wire [127:0] _add_map_x_29_all_sg_down;
  wire [127:0] _add_map_x_29_all_sg_right;
  wire [127:0] _add_map_x_29_all_sg_left;
  wire [7:0] _add_map_x_29_moto_org_near;
  wire [7:0] _add_map_x_29_moto_org_near1;
  wire [7:0] _add_map_x_29_moto_org_near2;
  wire [7:0] _add_map_x_29_moto_org_near3;
  wire [7:0] _add_map_x_29_moto_org;
  wire [1:0] _add_map_x_29_sg_up;
  wire [1:0] _add_map_x_29_sg_down;
  wire [1:0] _add_map_x_29_sg_left;
  wire [1:0] _add_map_x_29_sg_right;
  wire _add_map_x_29_wall_t_in;
  wire [7:0] _add_map_x_29_moto;
  wire [7:0] _add_map_x_29_up;
  wire [7:0] _add_map_x_29_right;
  wire [7:0] _add_map_x_29_down;
  wire [7:0] _add_map_x_29_left;
  wire [7:0] _add_map_x_29_start;
  wire [7:0] _add_map_x_29_goal;
  wire [7:0] _add_map_x_29_now;
  wire [7:0] _add_map_x_29_distance;
  wire [127:0] _add_map_x_29_end_wall;
  wire [127:0] _add_map_x_29_all_s_g;
  wire [127:0] _add_map_x_29_all_s_g_near;
  wire [7:0] _add_map_x_29_data_out;
  wire [7:0] _add_map_x_29_data_out_index;
  wire [7:0] _add_map_x_29_data_near;
  wire _add_map_x_29_wall_t_out;
  wire [7:0] _add_map_x_29_data_org;
  wire [7:0] _add_map_x_29_data_org_near;
  wire [1:0] _add_map_x_29_s_g;
  wire [1:0] _add_map_x_29_s_g_near;
  wire _add_map_x_29_add_exe;
  wire _add_map_x_29_p_reset;
  wire _add_map_x_29_m_clock;
  wire [127:0] _add_map_x_28_wall_end_in;
  wire [127:0] _add_map_x_28_all_sg_up;
  wire [127:0] _add_map_x_28_all_sg_down;
  wire [127:0] _add_map_x_28_all_sg_right;
  wire [127:0] _add_map_x_28_all_sg_left;
  wire [7:0] _add_map_x_28_moto_org_near;
  wire [7:0] _add_map_x_28_moto_org_near1;
  wire [7:0] _add_map_x_28_moto_org_near2;
  wire [7:0] _add_map_x_28_moto_org_near3;
  wire [7:0] _add_map_x_28_moto_org;
  wire [1:0] _add_map_x_28_sg_up;
  wire [1:0] _add_map_x_28_sg_down;
  wire [1:0] _add_map_x_28_sg_left;
  wire [1:0] _add_map_x_28_sg_right;
  wire _add_map_x_28_wall_t_in;
  wire [7:0] _add_map_x_28_moto;
  wire [7:0] _add_map_x_28_up;
  wire [7:0] _add_map_x_28_right;
  wire [7:0] _add_map_x_28_down;
  wire [7:0] _add_map_x_28_left;
  wire [7:0] _add_map_x_28_start;
  wire [7:0] _add_map_x_28_goal;
  wire [7:0] _add_map_x_28_now;
  wire [7:0] _add_map_x_28_distance;
  wire [127:0] _add_map_x_28_end_wall;
  wire [127:0] _add_map_x_28_all_s_g;
  wire [127:0] _add_map_x_28_all_s_g_near;
  wire [7:0] _add_map_x_28_data_out;
  wire [7:0] _add_map_x_28_data_out_index;
  wire [7:0] _add_map_x_28_data_near;
  wire _add_map_x_28_wall_t_out;
  wire [7:0] _add_map_x_28_data_org;
  wire [7:0] _add_map_x_28_data_org_near;
  wire [1:0] _add_map_x_28_s_g;
  wire [1:0] _add_map_x_28_s_g_near;
  wire _add_map_x_28_add_exe;
  wire _add_map_x_28_p_reset;
  wire _add_map_x_28_m_clock;
  wire [127:0] _add_map_x_27_wall_end_in;
  wire [127:0] _add_map_x_27_all_sg_up;
  wire [127:0] _add_map_x_27_all_sg_down;
  wire [127:0] _add_map_x_27_all_sg_right;
  wire [127:0] _add_map_x_27_all_sg_left;
  wire [7:0] _add_map_x_27_moto_org_near;
  wire [7:0] _add_map_x_27_moto_org_near1;
  wire [7:0] _add_map_x_27_moto_org_near2;
  wire [7:0] _add_map_x_27_moto_org_near3;
  wire [7:0] _add_map_x_27_moto_org;
  wire [1:0] _add_map_x_27_sg_up;
  wire [1:0] _add_map_x_27_sg_down;
  wire [1:0] _add_map_x_27_sg_left;
  wire [1:0] _add_map_x_27_sg_right;
  wire _add_map_x_27_wall_t_in;
  wire [7:0] _add_map_x_27_moto;
  wire [7:0] _add_map_x_27_up;
  wire [7:0] _add_map_x_27_right;
  wire [7:0] _add_map_x_27_down;
  wire [7:0] _add_map_x_27_left;
  wire [7:0] _add_map_x_27_start;
  wire [7:0] _add_map_x_27_goal;
  wire [7:0] _add_map_x_27_now;
  wire [7:0] _add_map_x_27_distance;
  wire [127:0] _add_map_x_27_end_wall;
  wire [127:0] _add_map_x_27_all_s_g;
  wire [127:0] _add_map_x_27_all_s_g_near;
  wire [7:0] _add_map_x_27_data_out;
  wire [7:0] _add_map_x_27_data_out_index;
  wire [7:0] _add_map_x_27_data_near;
  wire _add_map_x_27_wall_t_out;
  wire [7:0] _add_map_x_27_data_org;
  wire [7:0] _add_map_x_27_data_org_near;
  wire [1:0] _add_map_x_27_s_g;
  wire [1:0] _add_map_x_27_s_g_near;
  wire _add_map_x_27_add_exe;
  wire _add_map_x_27_p_reset;
  wire _add_map_x_27_m_clock;
  wire [127:0] _add_map_x_26_wall_end_in;
  wire [127:0] _add_map_x_26_all_sg_up;
  wire [127:0] _add_map_x_26_all_sg_down;
  wire [127:0] _add_map_x_26_all_sg_right;
  wire [127:0] _add_map_x_26_all_sg_left;
  wire [7:0] _add_map_x_26_moto_org_near;
  wire [7:0] _add_map_x_26_moto_org_near1;
  wire [7:0] _add_map_x_26_moto_org_near2;
  wire [7:0] _add_map_x_26_moto_org_near3;
  wire [7:0] _add_map_x_26_moto_org;
  wire [1:0] _add_map_x_26_sg_up;
  wire [1:0] _add_map_x_26_sg_down;
  wire [1:0] _add_map_x_26_sg_left;
  wire [1:0] _add_map_x_26_sg_right;
  wire _add_map_x_26_wall_t_in;
  wire [7:0] _add_map_x_26_moto;
  wire [7:0] _add_map_x_26_up;
  wire [7:0] _add_map_x_26_right;
  wire [7:0] _add_map_x_26_down;
  wire [7:0] _add_map_x_26_left;
  wire [7:0] _add_map_x_26_start;
  wire [7:0] _add_map_x_26_goal;
  wire [7:0] _add_map_x_26_now;
  wire [7:0] _add_map_x_26_distance;
  wire [127:0] _add_map_x_26_end_wall;
  wire [127:0] _add_map_x_26_all_s_g;
  wire [127:0] _add_map_x_26_all_s_g_near;
  wire [7:0] _add_map_x_26_data_out;
  wire [7:0] _add_map_x_26_data_out_index;
  wire [7:0] _add_map_x_26_data_near;
  wire _add_map_x_26_wall_t_out;
  wire [7:0] _add_map_x_26_data_org;
  wire [7:0] _add_map_x_26_data_org_near;
  wire [1:0] _add_map_x_26_s_g;
  wire [1:0] _add_map_x_26_s_g_near;
  wire _add_map_x_26_add_exe;
  wire _add_map_x_26_p_reset;
  wire _add_map_x_26_m_clock;
  wire [127:0] _add_map_x_25_wall_end_in;
  wire [127:0] _add_map_x_25_all_sg_up;
  wire [127:0] _add_map_x_25_all_sg_down;
  wire [127:0] _add_map_x_25_all_sg_right;
  wire [127:0] _add_map_x_25_all_sg_left;
  wire [7:0] _add_map_x_25_moto_org_near;
  wire [7:0] _add_map_x_25_moto_org_near1;
  wire [7:0] _add_map_x_25_moto_org_near2;
  wire [7:0] _add_map_x_25_moto_org_near3;
  wire [7:0] _add_map_x_25_moto_org;
  wire [1:0] _add_map_x_25_sg_up;
  wire [1:0] _add_map_x_25_sg_down;
  wire [1:0] _add_map_x_25_sg_left;
  wire [1:0] _add_map_x_25_sg_right;
  wire _add_map_x_25_wall_t_in;
  wire [7:0] _add_map_x_25_moto;
  wire [7:0] _add_map_x_25_up;
  wire [7:0] _add_map_x_25_right;
  wire [7:0] _add_map_x_25_down;
  wire [7:0] _add_map_x_25_left;
  wire [7:0] _add_map_x_25_start;
  wire [7:0] _add_map_x_25_goal;
  wire [7:0] _add_map_x_25_now;
  wire [7:0] _add_map_x_25_distance;
  wire [127:0] _add_map_x_25_end_wall;
  wire [127:0] _add_map_x_25_all_s_g;
  wire [127:0] _add_map_x_25_all_s_g_near;
  wire [7:0] _add_map_x_25_data_out;
  wire [7:0] _add_map_x_25_data_out_index;
  wire [7:0] _add_map_x_25_data_near;
  wire _add_map_x_25_wall_t_out;
  wire [7:0] _add_map_x_25_data_org;
  wire [7:0] _add_map_x_25_data_org_near;
  wire [1:0] _add_map_x_25_s_g;
  wire [1:0] _add_map_x_25_s_g_near;
  wire _add_map_x_25_add_exe;
  wire _add_map_x_25_p_reset;
  wire _add_map_x_25_m_clock;
  wire [127:0] _add_map_x_24_wall_end_in;
  wire [127:0] _add_map_x_24_all_sg_up;
  wire [127:0] _add_map_x_24_all_sg_down;
  wire [127:0] _add_map_x_24_all_sg_right;
  wire [127:0] _add_map_x_24_all_sg_left;
  wire [7:0] _add_map_x_24_moto_org_near;
  wire [7:0] _add_map_x_24_moto_org_near1;
  wire [7:0] _add_map_x_24_moto_org_near2;
  wire [7:0] _add_map_x_24_moto_org_near3;
  wire [7:0] _add_map_x_24_moto_org;
  wire [1:0] _add_map_x_24_sg_up;
  wire [1:0] _add_map_x_24_sg_down;
  wire [1:0] _add_map_x_24_sg_left;
  wire [1:0] _add_map_x_24_sg_right;
  wire _add_map_x_24_wall_t_in;
  wire [7:0] _add_map_x_24_moto;
  wire [7:0] _add_map_x_24_up;
  wire [7:0] _add_map_x_24_right;
  wire [7:0] _add_map_x_24_down;
  wire [7:0] _add_map_x_24_left;
  wire [7:0] _add_map_x_24_start;
  wire [7:0] _add_map_x_24_goal;
  wire [7:0] _add_map_x_24_now;
  wire [7:0] _add_map_x_24_distance;
  wire [127:0] _add_map_x_24_end_wall;
  wire [127:0] _add_map_x_24_all_s_g;
  wire [127:0] _add_map_x_24_all_s_g_near;
  wire [7:0] _add_map_x_24_data_out;
  wire [7:0] _add_map_x_24_data_out_index;
  wire [7:0] _add_map_x_24_data_near;
  wire _add_map_x_24_wall_t_out;
  wire [7:0] _add_map_x_24_data_org;
  wire [7:0] _add_map_x_24_data_org_near;
  wire [1:0] _add_map_x_24_s_g;
  wire [1:0] _add_map_x_24_s_g_near;
  wire _add_map_x_24_add_exe;
  wire _add_map_x_24_p_reset;
  wire _add_map_x_24_m_clock;
  wire [127:0] _add_map_x_23_wall_end_in;
  wire [127:0] _add_map_x_23_all_sg_up;
  wire [127:0] _add_map_x_23_all_sg_down;
  wire [127:0] _add_map_x_23_all_sg_right;
  wire [127:0] _add_map_x_23_all_sg_left;
  wire [7:0] _add_map_x_23_moto_org_near;
  wire [7:0] _add_map_x_23_moto_org_near1;
  wire [7:0] _add_map_x_23_moto_org_near2;
  wire [7:0] _add_map_x_23_moto_org_near3;
  wire [7:0] _add_map_x_23_moto_org;
  wire [1:0] _add_map_x_23_sg_up;
  wire [1:0] _add_map_x_23_sg_down;
  wire [1:0] _add_map_x_23_sg_left;
  wire [1:0] _add_map_x_23_sg_right;
  wire _add_map_x_23_wall_t_in;
  wire [7:0] _add_map_x_23_moto;
  wire [7:0] _add_map_x_23_up;
  wire [7:0] _add_map_x_23_right;
  wire [7:0] _add_map_x_23_down;
  wire [7:0] _add_map_x_23_left;
  wire [7:0] _add_map_x_23_start;
  wire [7:0] _add_map_x_23_goal;
  wire [7:0] _add_map_x_23_now;
  wire [7:0] _add_map_x_23_distance;
  wire [127:0] _add_map_x_23_end_wall;
  wire [127:0] _add_map_x_23_all_s_g;
  wire [127:0] _add_map_x_23_all_s_g_near;
  wire [7:0] _add_map_x_23_data_out;
  wire [7:0] _add_map_x_23_data_out_index;
  wire [7:0] _add_map_x_23_data_near;
  wire _add_map_x_23_wall_t_out;
  wire [7:0] _add_map_x_23_data_org;
  wire [7:0] _add_map_x_23_data_org_near;
  wire [1:0] _add_map_x_23_s_g;
  wire [1:0] _add_map_x_23_s_g_near;
  wire _add_map_x_23_add_exe;
  wire _add_map_x_23_p_reset;
  wire _add_map_x_23_m_clock;
  wire [127:0] _add_map_x_22_wall_end_in;
  wire [127:0] _add_map_x_22_all_sg_up;
  wire [127:0] _add_map_x_22_all_sg_down;
  wire [127:0] _add_map_x_22_all_sg_right;
  wire [127:0] _add_map_x_22_all_sg_left;
  wire [7:0] _add_map_x_22_moto_org_near;
  wire [7:0] _add_map_x_22_moto_org_near1;
  wire [7:0] _add_map_x_22_moto_org_near2;
  wire [7:0] _add_map_x_22_moto_org_near3;
  wire [7:0] _add_map_x_22_moto_org;
  wire [1:0] _add_map_x_22_sg_up;
  wire [1:0] _add_map_x_22_sg_down;
  wire [1:0] _add_map_x_22_sg_left;
  wire [1:0] _add_map_x_22_sg_right;
  wire _add_map_x_22_wall_t_in;
  wire [7:0] _add_map_x_22_moto;
  wire [7:0] _add_map_x_22_up;
  wire [7:0] _add_map_x_22_right;
  wire [7:0] _add_map_x_22_down;
  wire [7:0] _add_map_x_22_left;
  wire [7:0] _add_map_x_22_start;
  wire [7:0] _add_map_x_22_goal;
  wire [7:0] _add_map_x_22_now;
  wire [7:0] _add_map_x_22_distance;
  wire [127:0] _add_map_x_22_end_wall;
  wire [127:0] _add_map_x_22_all_s_g;
  wire [127:0] _add_map_x_22_all_s_g_near;
  wire [7:0] _add_map_x_22_data_out;
  wire [7:0] _add_map_x_22_data_out_index;
  wire [7:0] _add_map_x_22_data_near;
  wire _add_map_x_22_wall_t_out;
  wire [7:0] _add_map_x_22_data_org;
  wire [7:0] _add_map_x_22_data_org_near;
  wire [1:0] _add_map_x_22_s_g;
  wire [1:0] _add_map_x_22_s_g_near;
  wire _add_map_x_22_add_exe;
  wire _add_map_x_22_p_reset;
  wire _add_map_x_22_m_clock;
  wire [127:0] _add_map_x_21_wall_end_in;
  wire [127:0] _add_map_x_21_all_sg_up;
  wire [127:0] _add_map_x_21_all_sg_down;
  wire [127:0] _add_map_x_21_all_sg_right;
  wire [127:0] _add_map_x_21_all_sg_left;
  wire [7:0] _add_map_x_21_moto_org_near;
  wire [7:0] _add_map_x_21_moto_org_near1;
  wire [7:0] _add_map_x_21_moto_org_near2;
  wire [7:0] _add_map_x_21_moto_org_near3;
  wire [7:0] _add_map_x_21_moto_org;
  wire [1:0] _add_map_x_21_sg_up;
  wire [1:0] _add_map_x_21_sg_down;
  wire [1:0] _add_map_x_21_sg_left;
  wire [1:0] _add_map_x_21_sg_right;
  wire _add_map_x_21_wall_t_in;
  wire [7:0] _add_map_x_21_moto;
  wire [7:0] _add_map_x_21_up;
  wire [7:0] _add_map_x_21_right;
  wire [7:0] _add_map_x_21_down;
  wire [7:0] _add_map_x_21_left;
  wire [7:0] _add_map_x_21_start;
  wire [7:0] _add_map_x_21_goal;
  wire [7:0] _add_map_x_21_now;
  wire [7:0] _add_map_x_21_distance;
  wire [127:0] _add_map_x_21_end_wall;
  wire [127:0] _add_map_x_21_all_s_g;
  wire [127:0] _add_map_x_21_all_s_g_near;
  wire [7:0] _add_map_x_21_data_out;
  wire [7:0] _add_map_x_21_data_out_index;
  wire [7:0] _add_map_x_21_data_near;
  wire _add_map_x_21_wall_t_out;
  wire [7:0] _add_map_x_21_data_org;
  wire [7:0] _add_map_x_21_data_org_near;
  wire [1:0] _add_map_x_21_s_g;
  wire [1:0] _add_map_x_21_s_g_near;
  wire _add_map_x_21_add_exe;
  wire _add_map_x_21_p_reset;
  wire _add_map_x_21_m_clock;
  wire [127:0] _add_map_x_20_wall_end_in;
  wire [127:0] _add_map_x_20_all_sg_up;
  wire [127:0] _add_map_x_20_all_sg_down;
  wire [127:0] _add_map_x_20_all_sg_right;
  wire [127:0] _add_map_x_20_all_sg_left;
  wire [7:0] _add_map_x_20_moto_org_near;
  wire [7:0] _add_map_x_20_moto_org_near1;
  wire [7:0] _add_map_x_20_moto_org_near2;
  wire [7:0] _add_map_x_20_moto_org_near3;
  wire [7:0] _add_map_x_20_moto_org;
  wire [1:0] _add_map_x_20_sg_up;
  wire [1:0] _add_map_x_20_sg_down;
  wire [1:0] _add_map_x_20_sg_left;
  wire [1:0] _add_map_x_20_sg_right;
  wire _add_map_x_20_wall_t_in;
  wire [7:0] _add_map_x_20_moto;
  wire [7:0] _add_map_x_20_up;
  wire [7:0] _add_map_x_20_right;
  wire [7:0] _add_map_x_20_down;
  wire [7:0] _add_map_x_20_left;
  wire [7:0] _add_map_x_20_start;
  wire [7:0] _add_map_x_20_goal;
  wire [7:0] _add_map_x_20_now;
  wire [7:0] _add_map_x_20_distance;
  wire [127:0] _add_map_x_20_end_wall;
  wire [127:0] _add_map_x_20_all_s_g;
  wire [127:0] _add_map_x_20_all_s_g_near;
  wire [7:0] _add_map_x_20_data_out;
  wire [7:0] _add_map_x_20_data_out_index;
  wire [7:0] _add_map_x_20_data_near;
  wire _add_map_x_20_wall_t_out;
  wire [7:0] _add_map_x_20_data_org;
  wire [7:0] _add_map_x_20_data_org_near;
  wire [1:0] _add_map_x_20_s_g;
  wire [1:0] _add_map_x_20_s_g_near;
  wire _add_map_x_20_add_exe;
  wire _add_map_x_20_p_reset;
  wire _add_map_x_20_m_clock;
  wire [127:0] _add_map_x_19_wall_end_in;
  wire [127:0] _add_map_x_19_all_sg_up;
  wire [127:0] _add_map_x_19_all_sg_down;
  wire [127:0] _add_map_x_19_all_sg_right;
  wire [127:0] _add_map_x_19_all_sg_left;
  wire [7:0] _add_map_x_19_moto_org_near;
  wire [7:0] _add_map_x_19_moto_org_near1;
  wire [7:0] _add_map_x_19_moto_org_near2;
  wire [7:0] _add_map_x_19_moto_org_near3;
  wire [7:0] _add_map_x_19_moto_org;
  wire [1:0] _add_map_x_19_sg_up;
  wire [1:0] _add_map_x_19_sg_down;
  wire [1:0] _add_map_x_19_sg_left;
  wire [1:0] _add_map_x_19_sg_right;
  wire _add_map_x_19_wall_t_in;
  wire [7:0] _add_map_x_19_moto;
  wire [7:0] _add_map_x_19_up;
  wire [7:0] _add_map_x_19_right;
  wire [7:0] _add_map_x_19_down;
  wire [7:0] _add_map_x_19_left;
  wire [7:0] _add_map_x_19_start;
  wire [7:0] _add_map_x_19_goal;
  wire [7:0] _add_map_x_19_now;
  wire [7:0] _add_map_x_19_distance;
  wire [127:0] _add_map_x_19_end_wall;
  wire [127:0] _add_map_x_19_all_s_g;
  wire [127:0] _add_map_x_19_all_s_g_near;
  wire [7:0] _add_map_x_19_data_out;
  wire [7:0] _add_map_x_19_data_out_index;
  wire [7:0] _add_map_x_19_data_near;
  wire _add_map_x_19_wall_t_out;
  wire [7:0] _add_map_x_19_data_org;
  wire [7:0] _add_map_x_19_data_org_near;
  wire [1:0] _add_map_x_19_s_g;
  wire [1:0] _add_map_x_19_s_g_near;
  wire _add_map_x_19_add_exe;
  wire _add_map_x_19_p_reset;
  wire _add_map_x_19_m_clock;
  wire [127:0] _add_map_x_18_wall_end_in;
  wire [127:0] _add_map_x_18_all_sg_up;
  wire [127:0] _add_map_x_18_all_sg_down;
  wire [127:0] _add_map_x_18_all_sg_right;
  wire [127:0] _add_map_x_18_all_sg_left;
  wire [7:0] _add_map_x_18_moto_org_near;
  wire [7:0] _add_map_x_18_moto_org_near1;
  wire [7:0] _add_map_x_18_moto_org_near2;
  wire [7:0] _add_map_x_18_moto_org_near3;
  wire [7:0] _add_map_x_18_moto_org;
  wire [1:0] _add_map_x_18_sg_up;
  wire [1:0] _add_map_x_18_sg_down;
  wire [1:0] _add_map_x_18_sg_left;
  wire [1:0] _add_map_x_18_sg_right;
  wire _add_map_x_18_wall_t_in;
  wire [7:0] _add_map_x_18_moto;
  wire [7:0] _add_map_x_18_up;
  wire [7:0] _add_map_x_18_right;
  wire [7:0] _add_map_x_18_down;
  wire [7:0] _add_map_x_18_left;
  wire [7:0] _add_map_x_18_start;
  wire [7:0] _add_map_x_18_goal;
  wire [7:0] _add_map_x_18_now;
  wire [7:0] _add_map_x_18_distance;
  wire [127:0] _add_map_x_18_end_wall;
  wire [127:0] _add_map_x_18_all_s_g;
  wire [127:0] _add_map_x_18_all_s_g_near;
  wire [7:0] _add_map_x_18_data_out;
  wire [7:0] _add_map_x_18_data_out_index;
  wire [7:0] _add_map_x_18_data_near;
  wire _add_map_x_18_wall_t_out;
  wire [7:0] _add_map_x_18_data_org;
  wire [7:0] _add_map_x_18_data_org_near;
  wire [1:0] _add_map_x_18_s_g;
  wire [1:0] _add_map_x_18_s_g_near;
  wire _add_map_x_18_add_exe;
  wire _add_map_x_18_p_reset;
  wire _add_map_x_18_m_clock;
  wire [127:0] _add_map_x_17_wall_end_in;
  wire [127:0] _add_map_x_17_all_sg_up;
  wire [127:0] _add_map_x_17_all_sg_down;
  wire [127:0] _add_map_x_17_all_sg_right;
  wire [127:0] _add_map_x_17_all_sg_left;
  wire [7:0] _add_map_x_17_moto_org_near;
  wire [7:0] _add_map_x_17_moto_org_near1;
  wire [7:0] _add_map_x_17_moto_org_near2;
  wire [7:0] _add_map_x_17_moto_org_near3;
  wire [7:0] _add_map_x_17_moto_org;
  wire [1:0] _add_map_x_17_sg_up;
  wire [1:0] _add_map_x_17_sg_down;
  wire [1:0] _add_map_x_17_sg_left;
  wire [1:0] _add_map_x_17_sg_right;
  wire _add_map_x_17_wall_t_in;
  wire [7:0] _add_map_x_17_moto;
  wire [7:0] _add_map_x_17_up;
  wire [7:0] _add_map_x_17_right;
  wire [7:0] _add_map_x_17_down;
  wire [7:0] _add_map_x_17_left;
  wire [7:0] _add_map_x_17_start;
  wire [7:0] _add_map_x_17_goal;
  wire [7:0] _add_map_x_17_now;
  wire [7:0] _add_map_x_17_distance;
  wire [127:0] _add_map_x_17_end_wall;
  wire [127:0] _add_map_x_17_all_s_g;
  wire [127:0] _add_map_x_17_all_s_g_near;
  wire [7:0] _add_map_x_17_data_out;
  wire [7:0] _add_map_x_17_data_out_index;
  wire [7:0] _add_map_x_17_data_near;
  wire _add_map_x_17_wall_t_out;
  wire [7:0] _add_map_x_17_data_org;
  wire [7:0] _add_map_x_17_data_org_near;
  wire [1:0] _add_map_x_17_s_g;
  wire [1:0] _add_map_x_17_s_g_near;
  wire _add_map_x_17_add_exe;
  wire _add_map_x_17_p_reset;
  wire _add_map_x_17_m_clock;
  wire [127:0] _add_map_x_16_wall_end_in;
  wire [127:0] _add_map_x_16_all_sg_up;
  wire [127:0] _add_map_x_16_all_sg_down;
  wire [127:0] _add_map_x_16_all_sg_right;
  wire [127:0] _add_map_x_16_all_sg_left;
  wire [7:0] _add_map_x_16_moto_org_near;
  wire [7:0] _add_map_x_16_moto_org_near1;
  wire [7:0] _add_map_x_16_moto_org_near2;
  wire [7:0] _add_map_x_16_moto_org_near3;
  wire [7:0] _add_map_x_16_moto_org;
  wire [1:0] _add_map_x_16_sg_up;
  wire [1:0] _add_map_x_16_sg_down;
  wire [1:0] _add_map_x_16_sg_left;
  wire [1:0] _add_map_x_16_sg_right;
  wire _add_map_x_16_wall_t_in;
  wire [7:0] _add_map_x_16_moto;
  wire [7:0] _add_map_x_16_up;
  wire [7:0] _add_map_x_16_right;
  wire [7:0] _add_map_x_16_down;
  wire [7:0] _add_map_x_16_left;
  wire [7:0] _add_map_x_16_start;
  wire [7:0] _add_map_x_16_goal;
  wire [7:0] _add_map_x_16_now;
  wire [7:0] _add_map_x_16_distance;
  wire [127:0] _add_map_x_16_end_wall;
  wire [127:0] _add_map_x_16_all_s_g;
  wire [127:0] _add_map_x_16_all_s_g_near;
  wire [7:0] _add_map_x_16_data_out;
  wire [7:0] _add_map_x_16_data_out_index;
  wire [7:0] _add_map_x_16_data_near;
  wire _add_map_x_16_wall_t_out;
  wire [7:0] _add_map_x_16_data_org;
  wire [7:0] _add_map_x_16_data_org_near;
  wire [1:0] _add_map_x_16_s_g;
  wire [1:0] _add_map_x_16_s_g_near;
  wire _add_map_x_16_add_exe;
  wire _add_map_x_16_p_reset;
  wire _add_map_x_16_m_clock;
  wire [127:0] _add_map_x_15_wall_end_in;
  wire [127:0] _add_map_x_15_all_sg_up;
  wire [127:0] _add_map_x_15_all_sg_down;
  wire [127:0] _add_map_x_15_all_sg_right;
  wire [127:0] _add_map_x_15_all_sg_left;
  wire [7:0] _add_map_x_15_moto_org_near;
  wire [7:0] _add_map_x_15_moto_org_near1;
  wire [7:0] _add_map_x_15_moto_org_near2;
  wire [7:0] _add_map_x_15_moto_org_near3;
  wire [7:0] _add_map_x_15_moto_org;
  wire [1:0] _add_map_x_15_sg_up;
  wire [1:0] _add_map_x_15_sg_down;
  wire [1:0] _add_map_x_15_sg_left;
  wire [1:0] _add_map_x_15_sg_right;
  wire _add_map_x_15_wall_t_in;
  wire [7:0] _add_map_x_15_moto;
  wire [7:0] _add_map_x_15_up;
  wire [7:0] _add_map_x_15_right;
  wire [7:0] _add_map_x_15_down;
  wire [7:0] _add_map_x_15_left;
  wire [7:0] _add_map_x_15_start;
  wire [7:0] _add_map_x_15_goal;
  wire [7:0] _add_map_x_15_now;
  wire [7:0] _add_map_x_15_distance;
  wire [127:0] _add_map_x_15_end_wall;
  wire [127:0] _add_map_x_15_all_s_g;
  wire [127:0] _add_map_x_15_all_s_g_near;
  wire [7:0] _add_map_x_15_data_out;
  wire [7:0] _add_map_x_15_data_out_index;
  wire [7:0] _add_map_x_15_data_near;
  wire _add_map_x_15_wall_t_out;
  wire [7:0] _add_map_x_15_data_org;
  wire [7:0] _add_map_x_15_data_org_near;
  wire [1:0] _add_map_x_15_s_g;
  wire [1:0] _add_map_x_15_s_g_near;
  wire _add_map_x_15_add_exe;
  wire _add_map_x_15_p_reset;
  wire _add_map_x_15_m_clock;
  wire [127:0] _add_map_x_14_wall_end_in;
  wire [127:0] _add_map_x_14_all_sg_up;
  wire [127:0] _add_map_x_14_all_sg_down;
  wire [127:0] _add_map_x_14_all_sg_right;
  wire [127:0] _add_map_x_14_all_sg_left;
  wire [7:0] _add_map_x_14_moto_org_near;
  wire [7:0] _add_map_x_14_moto_org_near1;
  wire [7:0] _add_map_x_14_moto_org_near2;
  wire [7:0] _add_map_x_14_moto_org_near3;
  wire [7:0] _add_map_x_14_moto_org;
  wire [1:0] _add_map_x_14_sg_up;
  wire [1:0] _add_map_x_14_sg_down;
  wire [1:0] _add_map_x_14_sg_left;
  wire [1:0] _add_map_x_14_sg_right;
  wire _add_map_x_14_wall_t_in;
  wire [7:0] _add_map_x_14_moto;
  wire [7:0] _add_map_x_14_up;
  wire [7:0] _add_map_x_14_right;
  wire [7:0] _add_map_x_14_down;
  wire [7:0] _add_map_x_14_left;
  wire [7:0] _add_map_x_14_start;
  wire [7:0] _add_map_x_14_goal;
  wire [7:0] _add_map_x_14_now;
  wire [7:0] _add_map_x_14_distance;
  wire [127:0] _add_map_x_14_end_wall;
  wire [127:0] _add_map_x_14_all_s_g;
  wire [127:0] _add_map_x_14_all_s_g_near;
  wire [7:0] _add_map_x_14_data_out;
  wire [7:0] _add_map_x_14_data_out_index;
  wire [7:0] _add_map_x_14_data_near;
  wire _add_map_x_14_wall_t_out;
  wire [7:0] _add_map_x_14_data_org;
  wire [7:0] _add_map_x_14_data_org_near;
  wire [1:0] _add_map_x_14_s_g;
  wire [1:0] _add_map_x_14_s_g_near;
  wire _add_map_x_14_add_exe;
  wire _add_map_x_14_p_reset;
  wire _add_map_x_14_m_clock;
  wire [127:0] _add_map_x_13_wall_end_in;
  wire [127:0] _add_map_x_13_all_sg_up;
  wire [127:0] _add_map_x_13_all_sg_down;
  wire [127:0] _add_map_x_13_all_sg_right;
  wire [127:0] _add_map_x_13_all_sg_left;
  wire [7:0] _add_map_x_13_moto_org_near;
  wire [7:0] _add_map_x_13_moto_org_near1;
  wire [7:0] _add_map_x_13_moto_org_near2;
  wire [7:0] _add_map_x_13_moto_org_near3;
  wire [7:0] _add_map_x_13_moto_org;
  wire [1:0] _add_map_x_13_sg_up;
  wire [1:0] _add_map_x_13_sg_down;
  wire [1:0] _add_map_x_13_sg_left;
  wire [1:0] _add_map_x_13_sg_right;
  wire _add_map_x_13_wall_t_in;
  wire [7:0] _add_map_x_13_moto;
  wire [7:0] _add_map_x_13_up;
  wire [7:0] _add_map_x_13_right;
  wire [7:0] _add_map_x_13_down;
  wire [7:0] _add_map_x_13_left;
  wire [7:0] _add_map_x_13_start;
  wire [7:0] _add_map_x_13_goal;
  wire [7:0] _add_map_x_13_now;
  wire [7:0] _add_map_x_13_distance;
  wire [127:0] _add_map_x_13_end_wall;
  wire [127:0] _add_map_x_13_all_s_g;
  wire [127:0] _add_map_x_13_all_s_g_near;
  wire [7:0] _add_map_x_13_data_out;
  wire [7:0] _add_map_x_13_data_out_index;
  wire [7:0] _add_map_x_13_data_near;
  wire _add_map_x_13_wall_t_out;
  wire [7:0] _add_map_x_13_data_org;
  wire [7:0] _add_map_x_13_data_org_near;
  wire [1:0] _add_map_x_13_s_g;
  wire [1:0] _add_map_x_13_s_g_near;
  wire _add_map_x_13_add_exe;
  wire _add_map_x_13_p_reset;
  wire _add_map_x_13_m_clock;
  wire [127:0] _add_map_x_12_wall_end_in;
  wire [127:0] _add_map_x_12_all_sg_up;
  wire [127:0] _add_map_x_12_all_sg_down;
  wire [127:0] _add_map_x_12_all_sg_right;
  wire [127:0] _add_map_x_12_all_sg_left;
  wire [7:0] _add_map_x_12_moto_org_near;
  wire [7:0] _add_map_x_12_moto_org_near1;
  wire [7:0] _add_map_x_12_moto_org_near2;
  wire [7:0] _add_map_x_12_moto_org_near3;
  wire [7:0] _add_map_x_12_moto_org;
  wire [1:0] _add_map_x_12_sg_up;
  wire [1:0] _add_map_x_12_sg_down;
  wire [1:0] _add_map_x_12_sg_left;
  wire [1:0] _add_map_x_12_sg_right;
  wire _add_map_x_12_wall_t_in;
  wire [7:0] _add_map_x_12_moto;
  wire [7:0] _add_map_x_12_up;
  wire [7:0] _add_map_x_12_right;
  wire [7:0] _add_map_x_12_down;
  wire [7:0] _add_map_x_12_left;
  wire [7:0] _add_map_x_12_start;
  wire [7:0] _add_map_x_12_goal;
  wire [7:0] _add_map_x_12_now;
  wire [7:0] _add_map_x_12_distance;
  wire [127:0] _add_map_x_12_end_wall;
  wire [127:0] _add_map_x_12_all_s_g;
  wire [127:0] _add_map_x_12_all_s_g_near;
  wire [7:0] _add_map_x_12_data_out;
  wire [7:0] _add_map_x_12_data_out_index;
  wire [7:0] _add_map_x_12_data_near;
  wire _add_map_x_12_wall_t_out;
  wire [7:0] _add_map_x_12_data_org;
  wire [7:0] _add_map_x_12_data_org_near;
  wire [1:0] _add_map_x_12_s_g;
  wire [1:0] _add_map_x_12_s_g_near;
  wire _add_map_x_12_add_exe;
  wire _add_map_x_12_p_reset;
  wire _add_map_x_12_m_clock;
  wire [127:0] _add_map_x_11_wall_end_in;
  wire [127:0] _add_map_x_11_all_sg_up;
  wire [127:0] _add_map_x_11_all_sg_down;
  wire [127:0] _add_map_x_11_all_sg_right;
  wire [127:0] _add_map_x_11_all_sg_left;
  wire [7:0] _add_map_x_11_moto_org_near;
  wire [7:0] _add_map_x_11_moto_org_near1;
  wire [7:0] _add_map_x_11_moto_org_near2;
  wire [7:0] _add_map_x_11_moto_org_near3;
  wire [7:0] _add_map_x_11_moto_org;
  wire [1:0] _add_map_x_11_sg_up;
  wire [1:0] _add_map_x_11_sg_down;
  wire [1:0] _add_map_x_11_sg_left;
  wire [1:0] _add_map_x_11_sg_right;
  wire _add_map_x_11_wall_t_in;
  wire [7:0] _add_map_x_11_moto;
  wire [7:0] _add_map_x_11_up;
  wire [7:0] _add_map_x_11_right;
  wire [7:0] _add_map_x_11_down;
  wire [7:0] _add_map_x_11_left;
  wire [7:0] _add_map_x_11_start;
  wire [7:0] _add_map_x_11_goal;
  wire [7:0] _add_map_x_11_now;
  wire [7:0] _add_map_x_11_distance;
  wire [127:0] _add_map_x_11_end_wall;
  wire [127:0] _add_map_x_11_all_s_g;
  wire [127:0] _add_map_x_11_all_s_g_near;
  wire [7:0] _add_map_x_11_data_out;
  wire [7:0] _add_map_x_11_data_out_index;
  wire [7:0] _add_map_x_11_data_near;
  wire _add_map_x_11_wall_t_out;
  wire [7:0] _add_map_x_11_data_org;
  wire [7:0] _add_map_x_11_data_org_near;
  wire [1:0] _add_map_x_11_s_g;
  wire [1:0] _add_map_x_11_s_g_near;
  wire _add_map_x_11_add_exe;
  wire _add_map_x_11_p_reset;
  wire _add_map_x_11_m_clock;
  wire [127:0] _add_map_x_10_wall_end_in;
  wire [127:0] _add_map_x_10_all_sg_up;
  wire [127:0] _add_map_x_10_all_sg_down;
  wire [127:0] _add_map_x_10_all_sg_right;
  wire [127:0] _add_map_x_10_all_sg_left;
  wire [7:0] _add_map_x_10_moto_org_near;
  wire [7:0] _add_map_x_10_moto_org_near1;
  wire [7:0] _add_map_x_10_moto_org_near2;
  wire [7:0] _add_map_x_10_moto_org_near3;
  wire [7:0] _add_map_x_10_moto_org;
  wire [1:0] _add_map_x_10_sg_up;
  wire [1:0] _add_map_x_10_sg_down;
  wire [1:0] _add_map_x_10_sg_left;
  wire [1:0] _add_map_x_10_sg_right;
  wire _add_map_x_10_wall_t_in;
  wire [7:0] _add_map_x_10_moto;
  wire [7:0] _add_map_x_10_up;
  wire [7:0] _add_map_x_10_right;
  wire [7:0] _add_map_x_10_down;
  wire [7:0] _add_map_x_10_left;
  wire [7:0] _add_map_x_10_start;
  wire [7:0] _add_map_x_10_goal;
  wire [7:0] _add_map_x_10_now;
  wire [7:0] _add_map_x_10_distance;
  wire [127:0] _add_map_x_10_end_wall;
  wire [127:0] _add_map_x_10_all_s_g;
  wire [127:0] _add_map_x_10_all_s_g_near;
  wire [7:0] _add_map_x_10_data_out;
  wire [7:0] _add_map_x_10_data_out_index;
  wire [7:0] _add_map_x_10_data_near;
  wire _add_map_x_10_wall_t_out;
  wire [7:0] _add_map_x_10_data_org;
  wire [7:0] _add_map_x_10_data_org_near;
  wire [1:0] _add_map_x_10_s_g;
  wire [1:0] _add_map_x_10_s_g_near;
  wire _add_map_x_10_add_exe;
  wire _add_map_x_10_p_reset;
  wire _add_map_x_10_m_clock;
  wire [127:0] _add_map_x_9_wall_end_in;
  wire [127:0] _add_map_x_9_all_sg_up;
  wire [127:0] _add_map_x_9_all_sg_down;
  wire [127:0] _add_map_x_9_all_sg_right;
  wire [127:0] _add_map_x_9_all_sg_left;
  wire [7:0] _add_map_x_9_moto_org_near;
  wire [7:0] _add_map_x_9_moto_org_near1;
  wire [7:0] _add_map_x_9_moto_org_near2;
  wire [7:0] _add_map_x_9_moto_org_near3;
  wire [7:0] _add_map_x_9_moto_org;
  wire [1:0] _add_map_x_9_sg_up;
  wire [1:0] _add_map_x_9_sg_down;
  wire [1:0] _add_map_x_9_sg_left;
  wire [1:0] _add_map_x_9_sg_right;
  wire _add_map_x_9_wall_t_in;
  wire [7:0] _add_map_x_9_moto;
  wire [7:0] _add_map_x_9_up;
  wire [7:0] _add_map_x_9_right;
  wire [7:0] _add_map_x_9_down;
  wire [7:0] _add_map_x_9_left;
  wire [7:0] _add_map_x_9_start;
  wire [7:0] _add_map_x_9_goal;
  wire [7:0] _add_map_x_9_now;
  wire [7:0] _add_map_x_9_distance;
  wire [127:0] _add_map_x_9_end_wall;
  wire [127:0] _add_map_x_9_all_s_g;
  wire [127:0] _add_map_x_9_all_s_g_near;
  wire [7:0] _add_map_x_9_data_out;
  wire [7:0] _add_map_x_9_data_out_index;
  wire [7:0] _add_map_x_9_data_near;
  wire _add_map_x_9_wall_t_out;
  wire [7:0] _add_map_x_9_data_org;
  wire [7:0] _add_map_x_9_data_org_near;
  wire [1:0] _add_map_x_9_s_g;
  wire [1:0] _add_map_x_9_s_g_near;
  wire _add_map_x_9_add_exe;
  wire _add_map_x_9_p_reset;
  wire _add_map_x_9_m_clock;
  wire [127:0] _add_map_x_8_wall_end_in;
  wire [127:0] _add_map_x_8_all_sg_up;
  wire [127:0] _add_map_x_8_all_sg_down;
  wire [127:0] _add_map_x_8_all_sg_right;
  wire [127:0] _add_map_x_8_all_sg_left;
  wire [7:0] _add_map_x_8_moto_org_near;
  wire [7:0] _add_map_x_8_moto_org_near1;
  wire [7:0] _add_map_x_8_moto_org_near2;
  wire [7:0] _add_map_x_8_moto_org_near3;
  wire [7:0] _add_map_x_8_moto_org;
  wire [1:0] _add_map_x_8_sg_up;
  wire [1:0] _add_map_x_8_sg_down;
  wire [1:0] _add_map_x_8_sg_left;
  wire [1:0] _add_map_x_8_sg_right;
  wire _add_map_x_8_wall_t_in;
  wire [7:0] _add_map_x_8_moto;
  wire [7:0] _add_map_x_8_up;
  wire [7:0] _add_map_x_8_right;
  wire [7:0] _add_map_x_8_down;
  wire [7:0] _add_map_x_8_left;
  wire [7:0] _add_map_x_8_start;
  wire [7:0] _add_map_x_8_goal;
  wire [7:0] _add_map_x_8_now;
  wire [7:0] _add_map_x_8_distance;
  wire [127:0] _add_map_x_8_end_wall;
  wire [127:0] _add_map_x_8_all_s_g;
  wire [127:0] _add_map_x_8_all_s_g_near;
  wire [7:0] _add_map_x_8_data_out;
  wire [7:0] _add_map_x_8_data_out_index;
  wire [7:0] _add_map_x_8_data_near;
  wire _add_map_x_8_wall_t_out;
  wire [7:0] _add_map_x_8_data_org;
  wire [7:0] _add_map_x_8_data_org_near;
  wire [1:0] _add_map_x_8_s_g;
  wire [1:0] _add_map_x_8_s_g_near;
  wire _add_map_x_8_add_exe;
  wire _add_map_x_8_p_reset;
  wire _add_map_x_8_m_clock;
  wire [127:0] _add_map_x_7_wall_end_in;
  wire [127:0] _add_map_x_7_all_sg_up;
  wire [127:0] _add_map_x_7_all_sg_down;
  wire [127:0] _add_map_x_7_all_sg_right;
  wire [127:0] _add_map_x_7_all_sg_left;
  wire [7:0] _add_map_x_7_moto_org_near;
  wire [7:0] _add_map_x_7_moto_org_near1;
  wire [7:0] _add_map_x_7_moto_org_near2;
  wire [7:0] _add_map_x_7_moto_org_near3;
  wire [7:0] _add_map_x_7_moto_org;
  wire [1:0] _add_map_x_7_sg_up;
  wire [1:0] _add_map_x_7_sg_down;
  wire [1:0] _add_map_x_7_sg_left;
  wire [1:0] _add_map_x_7_sg_right;
  wire _add_map_x_7_wall_t_in;
  wire [7:0] _add_map_x_7_moto;
  wire [7:0] _add_map_x_7_up;
  wire [7:0] _add_map_x_7_right;
  wire [7:0] _add_map_x_7_down;
  wire [7:0] _add_map_x_7_left;
  wire [7:0] _add_map_x_7_start;
  wire [7:0] _add_map_x_7_goal;
  wire [7:0] _add_map_x_7_now;
  wire [7:0] _add_map_x_7_distance;
  wire [127:0] _add_map_x_7_end_wall;
  wire [127:0] _add_map_x_7_all_s_g;
  wire [127:0] _add_map_x_7_all_s_g_near;
  wire [7:0] _add_map_x_7_data_out;
  wire [7:0] _add_map_x_7_data_out_index;
  wire [7:0] _add_map_x_7_data_near;
  wire _add_map_x_7_wall_t_out;
  wire [7:0] _add_map_x_7_data_org;
  wire [7:0] _add_map_x_7_data_org_near;
  wire [1:0] _add_map_x_7_s_g;
  wire [1:0] _add_map_x_7_s_g_near;
  wire _add_map_x_7_add_exe;
  wire _add_map_x_7_p_reset;
  wire _add_map_x_7_m_clock;
  wire [127:0] _add_map_x_6_wall_end_in;
  wire [127:0] _add_map_x_6_all_sg_up;
  wire [127:0] _add_map_x_6_all_sg_down;
  wire [127:0] _add_map_x_6_all_sg_right;
  wire [127:0] _add_map_x_6_all_sg_left;
  wire [7:0] _add_map_x_6_moto_org_near;
  wire [7:0] _add_map_x_6_moto_org_near1;
  wire [7:0] _add_map_x_6_moto_org_near2;
  wire [7:0] _add_map_x_6_moto_org_near3;
  wire [7:0] _add_map_x_6_moto_org;
  wire [1:0] _add_map_x_6_sg_up;
  wire [1:0] _add_map_x_6_sg_down;
  wire [1:0] _add_map_x_6_sg_left;
  wire [1:0] _add_map_x_6_sg_right;
  wire _add_map_x_6_wall_t_in;
  wire [7:0] _add_map_x_6_moto;
  wire [7:0] _add_map_x_6_up;
  wire [7:0] _add_map_x_6_right;
  wire [7:0] _add_map_x_6_down;
  wire [7:0] _add_map_x_6_left;
  wire [7:0] _add_map_x_6_start;
  wire [7:0] _add_map_x_6_goal;
  wire [7:0] _add_map_x_6_now;
  wire [7:0] _add_map_x_6_distance;
  wire [127:0] _add_map_x_6_end_wall;
  wire [127:0] _add_map_x_6_all_s_g;
  wire [127:0] _add_map_x_6_all_s_g_near;
  wire [7:0] _add_map_x_6_data_out;
  wire [7:0] _add_map_x_6_data_out_index;
  wire [7:0] _add_map_x_6_data_near;
  wire _add_map_x_6_wall_t_out;
  wire [7:0] _add_map_x_6_data_org;
  wire [7:0] _add_map_x_6_data_org_near;
  wire [1:0] _add_map_x_6_s_g;
  wire [1:0] _add_map_x_6_s_g_near;
  wire _add_map_x_6_add_exe;
  wire _add_map_x_6_p_reset;
  wire _add_map_x_6_m_clock;
  wire [127:0] _add_map_x_5_wall_end_in;
  wire [127:0] _add_map_x_5_all_sg_up;
  wire [127:0] _add_map_x_5_all_sg_down;
  wire [127:0] _add_map_x_5_all_sg_right;
  wire [127:0] _add_map_x_5_all_sg_left;
  wire [7:0] _add_map_x_5_moto_org_near;
  wire [7:0] _add_map_x_5_moto_org_near1;
  wire [7:0] _add_map_x_5_moto_org_near2;
  wire [7:0] _add_map_x_5_moto_org_near3;
  wire [7:0] _add_map_x_5_moto_org;
  wire [1:0] _add_map_x_5_sg_up;
  wire [1:0] _add_map_x_5_sg_down;
  wire [1:0] _add_map_x_5_sg_left;
  wire [1:0] _add_map_x_5_sg_right;
  wire _add_map_x_5_wall_t_in;
  wire [7:0] _add_map_x_5_moto;
  wire [7:0] _add_map_x_5_up;
  wire [7:0] _add_map_x_5_right;
  wire [7:0] _add_map_x_5_down;
  wire [7:0] _add_map_x_5_left;
  wire [7:0] _add_map_x_5_start;
  wire [7:0] _add_map_x_5_goal;
  wire [7:0] _add_map_x_5_now;
  wire [7:0] _add_map_x_5_distance;
  wire [127:0] _add_map_x_5_end_wall;
  wire [127:0] _add_map_x_5_all_s_g;
  wire [127:0] _add_map_x_5_all_s_g_near;
  wire [7:0] _add_map_x_5_data_out;
  wire [7:0] _add_map_x_5_data_out_index;
  wire [7:0] _add_map_x_5_data_near;
  wire _add_map_x_5_wall_t_out;
  wire [7:0] _add_map_x_5_data_org;
  wire [7:0] _add_map_x_5_data_org_near;
  wire [1:0] _add_map_x_5_s_g;
  wire [1:0] _add_map_x_5_s_g_near;
  wire _add_map_x_5_add_exe;
  wire _add_map_x_5_p_reset;
  wire _add_map_x_5_m_clock;
  wire [127:0] _add_map_x_4_wall_end_in;
  wire [127:0] _add_map_x_4_all_sg_up;
  wire [127:0] _add_map_x_4_all_sg_down;
  wire [127:0] _add_map_x_4_all_sg_right;
  wire [127:0] _add_map_x_4_all_sg_left;
  wire [7:0] _add_map_x_4_moto_org_near;
  wire [7:0] _add_map_x_4_moto_org_near1;
  wire [7:0] _add_map_x_4_moto_org_near2;
  wire [7:0] _add_map_x_4_moto_org_near3;
  wire [7:0] _add_map_x_4_moto_org;
  wire [1:0] _add_map_x_4_sg_up;
  wire [1:0] _add_map_x_4_sg_down;
  wire [1:0] _add_map_x_4_sg_left;
  wire [1:0] _add_map_x_4_sg_right;
  wire _add_map_x_4_wall_t_in;
  wire [7:0] _add_map_x_4_moto;
  wire [7:0] _add_map_x_4_up;
  wire [7:0] _add_map_x_4_right;
  wire [7:0] _add_map_x_4_down;
  wire [7:0] _add_map_x_4_left;
  wire [7:0] _add_map_x_4_start;
  wire [7:0] _add_map_x_4_goal;
  wire [7:0] _add_map_x_4_now;
  wire [7:0] _add_map_x_4_distance;
  wire [127:0] _add_map_x_4_end_wall;
  wire [127:0] _add_map_x_4_all_s_g;
  wire [127:0] _add_map_x_4_all_s_g_near;
  wire [7:0] _add_map_x_4_data_out;
  wire [7:0] _add_map_x_4_data_out_index;
  wire [7:0] _add_map_x_4_data_near;
  wire _add_map_x_4_wall_t_out;
  wire [7:0] _add_map_x_4_data_org;
  wire [7:0] _add_map_x_4_data_org_near;
  wire [1:0] _add_map_x_4_s_g;
  wire [1:0] _add_map_x_4_s_g_near;
  wire _add_map_x_4_add_exe;
  wire _add_map_x_4_p_reset;
  wire _add_map_x_4_m_clock;
  wire [127:0] _add_map_x_3_wall_end_in;
  wire [127:0] _add_map_x_3_all_sg_up;
  wire [127:0] _add_map_x_3_all_sg_down;
  wire [127:0] _add_map_x_3_all_sg_right;
  wire [127:0] _add_map_x_3_all_sg_left;
  wire [7:0] _add_map_x_3_moto_org_near;
  wire [7:0] _add_map_x_3_moto_org_near1;
  wire [7:0] _add_map_x_3_moto_org_near2;
  wire [7:0] _add_map_x_3_moto_org_near3;
  wire [7:0] _add_map_x_3_moto_org;
  wire [1:0] _add_map_x_3_sg_up;
  wire [1:0] _add_map_x_3_sg_down;
  wire [1:0] _add_map_x_3_sg_left;
  wire [1:0] _add_map_x_3_sg_right;
  wire _add_map_x_3_wall_t_in;
  wire [7:0] _add_map_x_3_moto;
  wire [7:0] _add_map_x_3_up;
  wire [7:0] _add_map_x_3_right;
  wire [7:0] _add_map_x_3_down;
  wire [7:0] _add_map_x_3_left;
  wire [7:0] _add_map_x_3_start;
  wire [7:0] _add_map_x_3_goal;
  wire [7:0] _add_map_x_3_now;
  wire [7:0] _add_map_x_3_distance;
  wire [127:0] _add_map_x_3_end_wall;
  wire [127:0] _add_map_x_3_all_s_g;
  wire [127:0] _add_map_x_3_all_s_g_near;
  wire [7:0] _add_map_x_3_data_out;
  wire [7:0] _add_map_x_3_data_out_index;
  wire [7:0] _add_map_x_3_data_near;
  wire _add_map_x_3_wall_t_out;
  wire [7:0] _add_map_x_3_data_org;
  wire [7:0] _add_map_x_3_data_org_near;
  wire [1:0] _add_map_x_3_s_g;
  wire [1:0] _add_map_x_3_s_g_near;
  wire _add_map_x_3_add_exe;
  wire _add_map_x_3_p_reset;
  wire _add_map_x_3_m_clock;
  wire [127:0] _add_map_x_2_wall_end_in;
  wire [127:0] _add_map_x_2_all_sg_up;
  wire [127:0] _add_map_x_2_all_sg_down;
  wire [127:0] _add_map_x_2_all_sg_right;
  wire [127:0] _add_map_x_2_all_sg_left;
  wire [7:0] _add_map_x_2_moto_org_near;
  wire [7:0] _add_map_x_2_moto_org_near1;
  wire [7:0] _add_map_x_2_moto_org_near2;
  wire [7:0] _add_map_x_2_moto_org_near3;
  wire [7:0] _add_map_x_2_moto_org;
  wire [1:0] _add_map_x_2_sg_up;
  wire [1:0] _add_map_x_2_sg_down;
  wire [1:0] _add_map_x_2_sg_left;
  wire [1:0] _add_map_x_2_sg_right;
  wire _add_map_x_2_wall_t_in;
  wire [7:0] _add_map_x_2_moto;
  wire [7:0] _add_map_x_2_up;
  wire [7:0] _add_map_x_2_right;
  wire [7:0] _add_map_x_2_down;
  wire [7:0] _add_map_x_2_left;
  wire [7:0] _add_map_x_2_start;
  wire [7:0] _add_map_x_2_goal;
  wire [7:0] _add_map_x_2_now;
  wire [7:0] _add_map_x_2_distance;
  wire [127:0] _add_map_x_2_end_wall;
  wire [127:0] _add_map_x_2_all_s_g;
  wire [127:0] _add_map_x_2_all_s_g_near;
  wire [7:0] _add_map_x_2_data_out;
  wire [7:0] _add_map_x_2_data_out_index;
  wire [7:0] _add_map_x_2_data_near;
  wire _add_map_x_2_wall_t_out;
  wire [7:0] _add_map_x_2_data_org;
  wire [7:0] _add_map_x_2_data_org_near;
  wire [1:0] _add_map_x_2_s_g;
  wire [1:0] _add_map_x_2_s_g_near;
  wire _add_map_x_2_add_exe;
  wire _add_map_x_2_p_reset;
  wire _add_map_x_2_m_clock;
  wire [127:0] _add_map_x_1_wall_end_in;
  wire [127:0] _add_map_x_1_all_sg_up;
  wire [127:0] _add_map_x_1_all_sg_down;
  wire [127:0] _add_map_x_1_all_sg_right;
  wire [127:0] _add_map_x_1_all_sg_left;
  wire [7:0] _add_map_x_1_moto_org_near;
  wire [7:0] _add_map_x_1_moto_org_near1;
  wire [7:0] _add_map_x_1_moto_org_near2;
  wire [7:0] _add_map_x_1_moto_org_near3;
  wire [7:0] _add_map_x_1_moto_org;
  wire [1:0] _add_map_x_1_sg_up;
  wire [1:0] _add_map_x_1_sg_down;
  wire [1:0] _add_map_x_1_sg_left;
  wire [1:0] _add_map_x_1_sg_right;
  wire _add_map_x_1_wall_t_in;
  wire [7:0] _add_map_x_1_moto;
  wire [7:0] _add_map_x_1_up;
  wire [7:0] _add_map_x_1_right;
  wire [7:0] _add_map_x_1_down;
  wire [7:0] _add_map_x_1_left;
  wire [7:0] _add_map_x_1_start;
  wire [7:0] _add_map_x_1_goal;
  wire [7:0] _add_map_x_1_now;
  wire [7:0] _add_map_x_1_distance;
  wire [127:0] _add_map_x_1_end_wall;
  wire [127:0] _add_map_x_1_all_s_g;
  wire [127:0] _add_map_x_1_all_s_g_near;
  wire [7:0] _add_map_x_1_data_out;
  wire [7:0] _add_map_x_1_data_out_index;
  wire [7:0] _add_map_x_1_data_near;
  wire _add_map_x_1_wall_t_out;
  wire [7:0] _add_map_x_1_data_org;
  wire [7:0] _add_map_x_1_data_org_near;
  wire [1:0] _add_map_x_1_s_g;
  wire [1:0] _add_map_x_1_s_g_near;
  wire _add_map_x_1_add_exe;
  wire _add_map_x_1_p_reset;
  wire _add_map_x_1_m_clock;
  wire _net_0;
  wire _net_1;
  wire _net_2;
  wire _net_3;
add_map add_map_x (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_add_exe), .end_wall(_add_map_x_end_wall), .all_s_g(_add_map_x_all_s_g), .all_s_g_near(_add_map_x_all_s_g_near), .data_out(_add_map_x_data_out), .data_out_index(_add_map_x_data_out_index), .data_near(_add_map_x_data_near), .wall_t_out(_add_map_x_wall_t_out), .data_org(_add_map_x_data_org), .data_org_near(_add_map_x_data_org_near), .s_g(_add_map_x_s_g), .s_g_near(_add_map_x_s_g_near), .wall_end_in(_add_map_x_wall_end_in), .all_sg_up(_add_map_x_all_sg_up), .all_sg_down(_add_map_x_all_sg_down), .all_sg_right(_add_map_x_all_sg_right), .all_sg_left(_add_map_x_all_sg_left), .moto_org_near(_add_map_x_moto_org_near), .moto_org_near1(_add_map_x_moto_org_near1), .moto_org_near2(_add_map_x_moto_org_near2), .moto_org_near3(_add_map_x_moto_org_near3), .moto_org(_add_map_x_moto_org), .sg_up(_add_map_x_sg_up), .sg_down(_add_map_x_sg_down), .sg_left(_add_map_x_sg_left), .sg_right(_add_map_x_sg_right), .wall_t_in(_add_map_x_wall_t_in), .moto(_add_map_x_moto), .up(_add_map_x_up), .right(_add_map_x_right), .down(_add_map_x_down), .left(_add_map_x_left), .start(_add_map_x_start), .goal(_add_map_x_goal), .now(_add_map_x_now), .distance(_add_map_x_distance));
add_map add_map_x_41 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_41_add_exe), .end_wall(_add_map_x_41_end_wall), .all_s_g(_add_map_x_41_all_s_g), .all_s_g_near(_add_map_x_41_all_s_g_near), .data_out(_add_map_x_41_data_out), .data_out_index(_add_map_x_41_data_out_index), .data_near(_add_map_x_41_data_near), .wall_t_out(_add_map_x_41_wall_t_out), .data_org(_add_map_x_41_data_org), .data_org_near(_add_map_x_41_data_org_near), .s_g(_add_map_x_41_s_g), .s_g_near(_add_map_x_41_s_g_near), .wall_end_in(_add_map_x_41_wall_end_in), .all_sg_up(_add_map_x_41_all_sg_up), .all_sg_down(_add_map_x_41_all_sg_down), .all_sg_right(_add_map_x_41_all_sg_right), .all_sg_left(_add_map_x_41_all_sg_left), .moto_org_near(_add_map_x_41_moto_org_near), .moto_org_near1(_add_map_x_41_moto_org_near1), .moto_org_near2(_add_map_x_41_moto_org_near2), .moto_org_near3(_add_map_x_41_moto_org_near3), .moto_org(_add_map_x_41_moto_org), .sg_up(_add_map_x_41_sg_up), .sg_down(_add_map_x_41_sg_down), .sg_left(_add_map_x_41_sg_left), .sg_right(_add_map_x_41_sg_right), .wall_t_in(_add_map_x_41_wall_t_in), .moto(_add_map_x_41_moto), .up(_add_map_x_41_up), .right(_add_map_x_41_right), .down(_add_map_x_41_down), .left(_add_map_x_41_left), .start(_add_map_x_41_start), .goal(_add_map_x_41_goal), .now(_add_map_x_41_now), .distance(_add_map_x_41_distance));
add_map add_map_x_40 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_40_add_exe), .end_wall(_add_map_x_40_end_wall), .all_s_g(_add_map_x_40_all_s_g), .all_s_g_near(_add_map_x_40_all_s_g_near), .data_out(_add_map_x_40_data_out), .data_out_index(_add_map_x_40_data_out_index), .data_near(_add_map_x_40_data_near), .wall_t_out(_add_map_x_40_wall_t_out), .data_org(_add_map_x_40_data_org), .data_org_near(_add_map_x_40_data_org_near), .s_g(_add_map_x_40_s_g), .s_g_near(_add_map_x_40_s_g_near), .wall_end_in(_add_map_x_40_wall_end_in), .all_sg_up(_add_map_x_40_all_sg_up), .all_sg_down(_add_map_x_40_all_sg_down), .all_sg_right(_add_map_x_40_all_sg_right), .all_sg_left(_add_map_x_40_all_sg_left), .moto_org_near(_add_map_x_40_moto_org_near), .moto_org_near1(_add_map_x_40_moto_org_near1), .moto_org_near2(_add_map_x_40_moto_org_near2), .moto_org_near3(_add_map_x_40_moto_org_near3), .moto_org(_add_map_x_40_moto_org), .sg_up(_add_map_x_40_sg_up), .sg_down(_add_map_x_40_sg_down), .sg_left(_add_map_x_40_sg_left), .sg_right(_add_map_x_40_sg_right), .wall_t_in(_add_map_x_40_wall_t_in), .moto(_add_map_x_40_moto), .up(_add_map_x_40_up), .right(_add_map_x_40_right), .down(_add_map_x_40_down), .left(_add_map_x_40_left), .start(_add_map_x_40_start), .goal(_add_map_x_40_goal), .now(_add_map_x_40_now), .distance(_add_map_x_40_distance));
add_map add_map_x_39 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_39_add_exe), .end_wall(_add_map_x_39_end_wall), .all_s_g(_add_map_x_39_all_s_g), .all_s_g_near(_add_map_x_39_all_s_g_near), .data_out(_add_map_x_39_data_out), .data_out_index(_add_map_x_39_data_out_index), .data_near(_add_map_x_39_data_near), .wall_t_out(_add_map_x_39_wall_t_out), .data_org(_add_map_x_39_data_org), .data_org_near(_add_map_x_39_data_org_near), .s_g(_add_map_x_39_s_g), .s_g_near(_add_map_x_39_s_g_near), .wall_end_in(_add_map_x_39_wall_end_in), .all_sg_up(_add_map_x_39_all_sg_up), .all_sg_down(_add_map_x_39_all_sg_down), .all_sg_right(_add_map_x_39_all_sg_right), .all_sg_left(_add_map_x_39_all_sg_left), .moto_org_near(_add_map_x_39_moto_org_near), .moto_org_near1(_add_map_x_39_moto_org_near1), .moto_org_near2(_add_map_x_39_moto_org_near2), .moto_org_near3(_add_map_x_39_moto_org_near3), .moto_org(_add_map_x_39_moto_org), .sg_up(_add_map_x_39_sg_up), .sg_down(_add_map_x_39_sg_down), .sg_left(_add_map_x_39_sg_left), .sg_right(_add_map_x_39_sg_right), .wall_t_in(_add_map_x_39_wall_t_in), .moto(_add_map_x_39_moto), .up(_add_map_x_39_up), .right(_add_map_x_39_right), .down(_add_map_x_39_down), .left(_add_map_x_39_left), .start(_add_map_x_39_start), .goal(_add_map_x_39_goal), .now(_add_map_x_39_now), .distance(_add_map_x_39_distance));
add_map add_map_x_38 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_38_add_exe), .end_wall(_add_map_x_38_end_wall), .all_s_g(_add_map_x_38_all_s_g), .all_s_g_near(_add_map_x_38_all_s_g_near), .data_out(_add_map_x_38_data_out), .data_out_index(_add_map_x_38_data_out_index), .data_near(_add_map_x_38_data_near), .wall_t_out(_add_map_x_38_wall_t_out), .data_org(_add_map_x_38_data_org), .data_org_near(_add_map_x_38_data_org_near), .s_g(_add_map_x_38_s_g), .s_g_near(_add_map_x_38_s_g_near), .wall_end_in(_add_map_x_38_wall_end_in), .all_sg_up(_add_map_x_38_all_sg_up), .all_sg_down(_add_map_x_38_all_sg_down), .all_sg_right(_add_map_x_38_all_sg_right), .all_sg_left(_add_map_x_38_all_sg_left), .moto_org_near(_add_map_x_38_moto_org_near), .moto_org_near1(_add_map_x_38_moto_org_near1), .moto_org_near2(_add_map_x_38_moto_org_near2), .moto_org_near3(_add_map_x_38_moto_org_near3), .moto_org(_add_map_x_38_moto_org), .sg_up(_add_map_x_38_sg_up), .sg_down(_add_map_x_38_sg_down), .sg_left(_add_map_x_38_sg_left), .sg_right(_add_map_x_38_sg_right), .wall_t_in(_add_map_x_38_wall_t_in), .moto(_add_map_x_38_moto), .up(_add_map_x_38_up), .right(_add_map_x_38_right), .down(_add_map_x_38_down), .left(_add_map_x_38_left), .start(_add_map_x_38_start), .goal(_add_map_x_38_goal), .now(_add_map_x_38_now), .distance(_add_map_x_38_distance));
add_map add_map_x_37 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_37_add_exe), .end_wall(_add_map_x_37_end_wall), .all_s_g(_add_map_x_37_all_s_g), .all_s_g_near(_add_map_x_37_all_s_g_near), .data_out(_add_map_x_37_data_out), .data_out_index(_add_map_x_37_data_out_index), .data_near(_add_map_x_37_data_near), .wall_t_out(_add_map_x_37_wall_t_out), .data_org(_add_map_x_37_data_org), .data_org_near(_add_map_x_37_data_org_near), .s_g(_add_map_x_37_s_g), .s_g_near(_add_map_x_37_s_g_near), .wall_end_in(_add_map_x_37_wall_end_in), .all_sg_up(_add_map_x_37_all_sg_up), .all_sg_down(_add_map_x_37_all_sg_down), .all_sg_right(_add_map_x_37_all_sg_right), .all_sg_left(_add_map_x_37_all_sg_left), .moto_org_near(_add_map_x_37_moto_org_near), .moto_org_near1(_add_map_x_37_moto_org_near1), .moto_org_near2(_add_map_x_37_moto_org_near2), .moto_org_near3(_add_map_x_37_moto_org_near3), .moto_org(_add_map_x_37_moto_org), .sg_up(_add_map_x_37_sg_up), .sg_down(_add_map_x_37_sg_down), .sg_left(_add_map_x_37_sg_left), .sg_right(_add_map_x_37_sg_right), .wall_t_in(_add_map_x_37_wall_t_in), .moto(_add_map_x_37_moto), .up(_add_map_x_37_up), .right(_add_map_x_37_right), .down(_add_map_x_37_down), .left(_add_map_x_37_left), .start(_add_map_x_37_start), .goal(_add_map_x_37_goal), .now(_add_map_x_37_now), .distance(_add_map_x_37_distance));
add_map add_map_x_36 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_36_add_exe), .end_wall(_add_map_x_36_end_wall), .all_s_g(_add_map_x_36_all_s_g), .all_s_g_near(_add_map_x_36_all_s_g_near), .data_out(_add_map_x_36_data_out), .data_out_index(_add_map_x_36_data_out_index), .data_near(_add_map_x_36_data_near), .wall_t_out(_add_map_x_36_wall_t_out), .data_org(_add_map_x_36_data_org), .data_org_near(_add_map_x_36_data_org_near), .s_g(_add_map_x_36_s_g), .s_g_near(_add_map_x_36_s_g_near), .wall_end_in(_add_map_x_36_wall_end_in), .all_sg_up(_add_map_x_36_all_sg_up), .all_sg_down(_add_map_x_36_all_sg_down), .all_sg_right(_add_map_x_36_all_sg_right), .all_sg_left(_add_map_x_36_all_sg_left), .moto_org_near(_add_map_x_36_moto_org_near), .moto_org_near1(_add_map_x_36_moto_org_near1), .moto_org_near2(_add_map_x_36_moto_org_near2), .moto_org_near3(_add_map_x_36_moto_org_near3), .moto_org(_add_map_x_36_moto_org), .sg_up(_add_map_x_36_sg_up), .sg_down(_add_map_x_36_sg_down), .sg_left(_add_map_x_36_sg_left), .sg_right(_add_map_x_36_sg_right), .wall_t_in(_add_map_x_36_wall_t_in), .moto(_add_map_x_36_moto), .up(_add_map_x_36_up), .right(_add_map_x_36_right), .down(_add_map_x_36_down), .left(_add_map_x_36_left), .start(_add_map_x_36_start), .goal(_add_map_x_36_goal), .now(_add_map_x_36_now), .distance(_add_map_x_36_distance));
add_map add_map_x_35 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_35_add_exe), .end_wall(_add_map_x_35_end_wall), .all_s_g(_add_map_x_35_all_s_g), .all_s_g_near(_add_map_x_35_all_s_g_near), .data_out(_add_map_x_35_data_out), .data_out_index(_add_map_x_35_data_out_index), .data_near(_add_map_x_35_data_near), .wall_t_out(_add_map_x_35_wall_t_out), .data_org(_add_map_x_35_data_org), .data_org_near(_add_map_x_35_data_org_near), .s_g(_add_map_x_35_s_g), .s_g_near(_add_map_x_35_s_g_near), .wall_end_in(_add_map_x_35_wall_end_in), .all_sg_up(_add_map_x_35_all_sg_up), .all_sg_down(_add_map_x_35_all_sg_down), .all_sg_right(_add_map_x_35_all_sg_right), .all_sg_left(_add_map_x_35_all_sg_left), .moto_org_near(_add_map_x_35_moto_org_near), .moto_org_near1(_add_map_x_35_moto_org_near1), .moto_org_near2(_add_map_x_35_moto_org_near2), .moto_org_near3(_add_map_x_35_moto_org_near3), .moto_org(_add_map_x_35_moto_org), .sg_up(_add_map_x_35_sg_up), .sg_down(_add_map_x_35_sg_down), .sg_left(_add_map_x_35_sg_left), .sg_right(_add_map_x_35_sg_right), .wall_t_in(_add_map_x_35_wall_t_in), .moto(_add_map_x_35_moto), .up(_add_map_x_35_up), .right(_add_map_x_35_right), .down(_add_map_x_35_down), .left(_add_map_x_35_left), .start(_add_map_x_35_start), .goal(_add_map_x_35_goal), .now(_add_map_x_35_now), .distance(_add_map_x_35_distance));
add_map add_map_x_34 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_34_add_exe), .end_wall(_add_map_x_34_end_wall), .all_s_g(_add_map_x_34_all_s_g), .all_s_g_near(_add_map_x_34_all_s_g_near), .data_out(_add_map_x_34_data_out), .data_out_index(_add_map_x_34_data_out_index), .data_near(_add_map_x_34_data_near), .wall_t_out(_add_map_x_34_wall_t_out), .data_org(_add_map_x_34_data_org), .data_org_near(_add_map_x_34_data_org_near), .s_g(_add_map_x_34_s_g), .s_g_near(_add_map_x_34_s_g_near), .wall_end_in(_add_map_x_34_wall_end_in), .all_sg_up(_add_map_x_34_all_sg_up), .all_sg_down(_add_map_x_34_all_sg_down), .all_sg_right(_add_map_x_34_all_sg_right), .all_sg_left(_add_map_x_34_all_sg_left), .moto_org_near(_add_map_x_34_moto_org_near), .moto_org_near1(_add_map_x_34_moto_org_near1), .moto_org_near2(_add_map_x_34_moto_org_near2), .moto_org_near3(_add_map_x_34_moto_org_near3), .moto_org(_add_map_x_34_moto_org), .sg_up(_add_map_x_34_sg_up), .sg_down(_add_map_x_34_sg_down), .sg_left(_add_map_x_34_sg_left), .sg_right(_add_map_x_34_sg_right), .wall_t_in(_add_map_x_34_wall_t_in), .moto(_add_map_x_34_moto), .up(_add_map_x_34_up), .right(_add_map_x_34_right), .down(_add_map_x_34_down), .left(_add_map_x_34_left), .start(_add_map_x_34_start), .goal(_add_map_x_34_goal), .now(_add_map_x_34_now), .distance(_add_map_x_34_distance));
add_map add_map_x_33 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_33_add_exe), .end_wall(_add_map_x_33_end_wall), .all_s_g(_add_map_x_33_all_s_g), .all_s_g_near(_add_map_x_33_all_s_g_near), .data_out(_add_map_x_33_data_out), .data_out_index(_add_map_x_33_data_out_index), .data_near(_add_map_x_33_data_near), .wall_t_out(_add_map_x_33_wall_t_out), .data_org(_add_map_x_33_data_org), .data_org_near(_add_map_x_33_data_org_near), .s_g(_add_map_x_33_s_g), .s_g_near(_add_map_x_33_s_g_near), .wall_end_in(_add_map_x_33_wall_end_in), .all_sg_up(_add_map_x_33_all_sg_up), .all_sg_down(_add_map_x_33_all_sg_down), .all_sg_right(_add_map_x_33_all_sg_right), .all_sg_left(_add_map_x_33_all_sg_left), .moto_org_near(_add_map_x_33_moto_org_near), .moto_org_near1(_add_map_x_33_moto_org_near1), .moto_org_near2(_add_map_x_33_moto_org_near2), .moto_org_near3(_add_map_x_33_moto_org_near3), .moto_org(_add_map_x_33_moto_org), .sg_up(_add_map_x_33_sg_up), .sg_down(_add_map_x_33_sg_down), .sg_left(_add_map_x_33_sg_left), .sg_right(_add_map_x_33_sg_right), .wall_t_in(_add_map_x_33_wall_t_in), .moto(_add_map_x_33_moto), .up(_add_map_x_33_up), .right(_add_map_x_33_right), .down(_add_map_x_33_down), .left(_add_map_x_33_left), .start(_add_map_x_33_start), .goal(_add_map_x_33_goal), .now(_add_map_x_33_now), .distance(_add_map_x_33_distance));
add_map add_map_x_32 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_32_add_exe), .end_wall(_add_map_x_32_end_wall), .all_s_g(_add_map_x_32_all_s_g), .all_s_g_near(_add_map_x_32_all_s_g_near), .data_out(_add_map_x_32_data_out), .data_out_index(_add_map_x_32_data_out_index), .data_near(_add_map_x_32_data_near), .wall_t_out(_add_map_x_32_wall_t_out), .data_org(_add_map_x_32_data_org), .data_org_near(_add_map_x_32_data_org_near), .s_g(_add_map_x_32_s_g), .s_g_near(_add_map_x_32_s_g_near), .wall_end_in(_add_map_x_32_wall_end_in), .all_sg_up(_add_map_x_32_all_sg_up), .all_sg_down(_add_map_x_32_all_sg_down), .all_sg_right(_add_map_x_32_all_sg_right), .all_sg_left(_add_map_x_32_all_sg_left), .moto_org_near(_add_map_x_32_moto_org_near), .moto_org_near1(_add_map_x_32_moto_org_near1), .moto_org_near2(_add_map_x_32_moto_org_near2), .moto_org_near3(_add_map_x_32_moto_org_near3), .moto_org(_add_map_x_32_moto_org), .sg_up(_add_map_x_32_sg_up), .sg_down(_add_map_x_32_sg_down), .sg_left(_add_map_x_32_sg_left), .sg_right(_add_map_x_32_sg_right), .wall_t_in(_add_map_x_32_wall_t_in), .moto(_add_map_x_32_moto), .up(_add_map_x_32_up), .right(_add_map_x_32_right), .down(_add_map_x_32_down), .left(_add_map_x_32_left), .start(_add_map_x_32_start), .goal(_add_map_x_32_goal), .now(_add_map_x_32_now), .distance(_add_map_x_32_distance));
add_map add_map_x_31 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_31_add_exe), .end_wall(_add_map_x_31_end_wall), .all_s_g(_add_map_x_31_all_s_g), .all_s_g_near(_add_map_x_31_all_s_g_near), .data_out(_add_map_x_31_data_out), .data_out_index(_add_map_x_31_data_out_index), .data_near(_add_map_x_31_data_near), .wall_t_out(_add_map_x_31_wall_t_out), .data_org(_add_map_x_31_data_org), .data_org_near(_add_map_x_31_data_org_near), .s_g(_add_map_x_31_s_g), .s_g_near(_add_map_x_31_s_g_near), .wall_end_in(_add_map_x_31_wall_end_in), .all_sg_up(_add_map_x_31_all_sg_up), .all_sg_down(_add_map_x_31_all_sg_down), .all_sg_right(_add_map_x_31_all_sg_right), .all_sg_left(_add_map_x_31_all_sg_left), .moto_org_near(_add_map_x_31_moto_org_near), .moto_org_near1(_add_map_x_31_moto_org_near1), .moto_org_near2(_add_map_x_31_moto_org_near2), .moto_org_near3(_add_map_x_31_moto_org_near3), .moto_org(_add_map_x_31_moto_org), .sg_up(_add_map_x_31_sg_up), .sg_down(_add_map_x_31_sg_down), .sg_left(_add_map_x_31_sg_left), .sg_right(_add_map_x_31_sg_right), .wall_t_in(_add_map_x_31_wall_t_in), .moto(_add_map_x_31_moto), .up(_add_map_x_31_up), .right(_add_map_x_31_right), .down(_add_map_x_31_down), .left(_add_map_x_31_left), .start(_add_map_x_31_start), .goal(_add_map_x_31_goal), .now(_add_map_x_31_now), .distance(_add_map_x_31_distance));
add_map add_map_x_30 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_30_add_exe), .end_wall(_add_map_x_30_end_wall), .all_s_g(_add_map_x_30_all_s_g), .all_s_g_near(_add_map_x_30_all_s_g_near), .data_out(_add_map_x_30_data_out), .data_out_index(_add_map_x_30_data_out_index), .data_near(_add_map_x_30_data_near), .wall_t_out(_add_map_x_30_wall_t_out), .data_org(_add_map_x_30_data_org), .data_org_near(_add_map_x_30_data_org_near), .s_g(_add_map_x_30_s_g), .s_g_near(_add_map_x_30_s_g_near), .wall_end_in(_add_map_x_30_wall_end_in), .all_sg_up(_add_map_x_30_all_sg_up), .all_sg_down(_add_map_x_30_all_sg_down), .all_sg_right(_add_map_x_30_all_sg_right), .all_sg_left(_add_map_x_30_all_sg_left), .moto_org_near(_add_map_x_30_moto_org_near), .moto_org_near1(_add_map_x_30_moto_org_near1), .moto_org_near2(_add_map_x_30_moto_org_near2), .moto_org_near3(_add_map_x_30_moto_org_near3), .moto_org(_add_map_x_30_moto_org), .sg_up(_add_map_x_30_sg_up), .sg_down(_add_map_x_30_sg_down), .sg_left(_add_map_x_30_sg_left), .sg_right(_add_map_x_30_sg_right), .wall_t_in(_add_map_x_30_wall_t_in), .moto(_add_map_x_30_moto), .up(_add_map_x_30_up), .right(_add_map_x_30_right), .down(_add_map_x_30_down), .left(_add_map_x_30_left), .start(_add_map_x_30_start), .goal(_add_map_x_30_goal), .now(_add_map_x_30_now), .distance(_add_map_x_30_distance));
add_map add_map_x_29 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_29_add_exe), .end_wall(_add_map_x_29_end_wall), .all_s_g(_add_map_x_29_all_s_g), .all_s_g_near(_add_map_x_29_all_s_g_near), .data_out(_add_map_x_29_data_out), .data_out_index(_add_map_x_29_data_out_index), .data_near(_add_map_x_29_data_near), .wall_t_out(_add_map_x_29_wall_t_out), .data_org(_add_map_x_29_data_org), .data_org_near(_add_map_x_29_data_org_near), .s_g(_add_map_x_29_s_g), .s_g_near(_add_map_x_29_s_g_near), .wall_end_in(_add_map_x_29_wall_end_in), .all_sg_up(_add_map_x_29_all_sg_up), .all_sg_down(_add_map_x_29_all_sg_down), .all_sg_right(_add_map_x_29_all_sg_right), .all_sg_left(_add_map_x_29_all_sg_left), .moto_org_near(_add_map_x_29_moto_org_near), .moto_org_near1(_add_map_x_29_moto_org_near1), .moto_org_near2(_add_map_x_29_moto_org_near2), .moto_org_near3(_add_map_x_29_moto_org_near3), .moto_org(_add_map_x_29_moto_org), .sg_up(_add_map_x_29_sg_up), .sg_down(_add_map_x_29_sg_down), .sg_left(_add_map_x_29_sg_left), .sg_right(_add_map_x_29_sg_right), .wall_t_in(_add_map_x_29_wall_t_in), .moto(_add_map_x_29_moto), .up(_add_map_x_29_up), .right(_add_map_x_29_right), .down(_add_map_x_29_down), .left(_add_map_x_29_left), .start(_add_map_x_29_start), .goal(_add_map_x_29_goal), .now(_add_map_x_29_now), .distance(_add_map_x_29_distance));
add_map add_map_x_28 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_28_add_exe), .end_wall(_add_map_x_28_end_wall), .all_s_g(_add_map_x_28_all_s_g), .all_s_g_near(_add_map_x_28_all_s_g_near), .data_out(_add_map_x_28_data_out), .data_out_index(_add_map_x_28_data_out_index), .data_near(_add_map_x_28_data_near), .wall_t_out(_add_map_x_28_wall_t_out), .data_org(_add_map_x_28_data_org), .data_org_near(_add_map_x_28_data_org_near), .s_g(_add_map_x_28_s_g), .s_g_near(_add_map_x_28_s_g_near), .wall_end_in(_add_map_x_28_wall_end_in), .all_sg_up(_add_map_x_28_all_sg_up), .all_sg_down(_add_map_x_28_all_sg_down), .all_sg_right(_add_map_x_28_all_sg_right), .all_sg_left(_add_map_x_28_all_sg_left), .moto_org_near(_add_map_x_28_moto_org_near), .moto_org_near1(_add_map_x_28_moto_org_near1), .moto_org_near2(_add_map_x_28_moto_org_near2), .moto_org_near3(_add_map_x_28_moto_org_near3), .moto_org(_add_map_x_28_moto_org), .sg_up(_add_map_x_28_sg_up), .sg_down(_add_map_x_28_sg_down), .sg_left(_add_map_x_28_sg_left), .sg_right(_add_map_x_28_sg_right), .wall_t_in(_add_map_x_28_wall_t_in), .moto(_add_map_x_28_moto), .up(_add_map_x_28_up), .right(_add_map_x_28_right), .down(_add_map_x_28_down), .left(_add_map_x_28_left), .start(_add_map_x_28_start), .goal(_add_map_x_28_goal), .now(_add_map_x_28_now), .distance(_add_map_x_28_distance));
add_map add_map_x_27 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_27_add_exe), .end_wall(_add_map_x_27_end_wall), .all_s_g(_add_map_x_27_all_s_g), .all_s_g_near(_add_map_x_27_all_s_g_near), .data_out(_add_map_x_27_data_out), .data_out_index(_add_map_x_27_data_out_index), .data_near(_add_map_x_27_data_near), .wall_t_out(_add_map_x_27_wall_t_out), .data_org(_add_map_x_27_data_org), .data_org_near(_add_map_x_27_data_org_near), .s_g(_add_map_x_27_s_g), .s_g_near(_add_map_x_27_s_g_near), .wall_end_in(_add_map_x_27_wall_end_in), .all_sg_up(_add_map_x_27_all_sg_up), .all_sg_down(_add_map_x_27_all_sg_down), .all_sg_right(_add_map_x_27_all_sg_right), .all_sg_left(_add_map_x_27_all_sg_left), .moto_org_near(_add_map_x_27_moto_org_near), .moto_org_near1(_add_map_x_27_moto_org_near1), .moto_org_near2(_add_map_x_27_moto_org_near2), .moto_org_near3(_add_map_x_27_moto_org_near3), .moto_org(_add_map_x_27_moto_org), .sg_up(_add_map_x_27_sg_up), .sg_down(_add_map_x_27_sg_down), .sg_left(_add_map_x_27_sg_left), .sg_right(_add_map_x_27_sg_right), .wall_t_in(_add_map_x_27_wall_t_in), .moto(_add_map_x_27_moto), .up(_add_map_x_27_up), .right(_add_map_x_27_right), .down(_add_map_x_27_down), .left(_add_map_x_27_left), .start(_add_map_x_27_start), .goal(_add_map_x_27_goal), .now(_add_map_x_27_now), .distance(_add_map_x_27_distance));
add_map add_map_x_26 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_26_add_exe), .end_wall(_add_map_x_26_end_wall), .all_s_g(_add_map_x_26_all_s_g), .all_s_g_near(_add_map_x_26_all_s_g_near), .data_out(_add_map_x_26_data_out), .data_out_index(_add_map_x_26_data_out_index), .data_near(_add_map_x_26_data_near), .wall_t_out(_add_map_x_26_wall_t_out), .data_org(_add_map_x_26_data_org), .data_org_near(_add_map_x_26_data_org_near), .s_g(_add_map_x_26_s_g), .s_g_near(_add_map_x_26_s_g_near), .wall_end_in(_add_map_x_26_wall_end_in), .all_sg_up(_add_map_x_26_all_sg_up), .all_sg_down(_add_map_x_26_all_sg_down), .all_sg_right(_add_map_x_26_all_sg_right), .all_sg_left(_add_map_x_26_all_sg_left), .moto_org_near(_add_map_x_26_moto_org_near), .moto_org_near1(_add_map_x_26_moto_org_near1), .moto_org_near2(_add_map_x_26_moto_org_near2), .moto_org_near3(_add_map_x_26_moto_org_near3), .moto_org(_add_map_x_26_moto_org), .sg_up(_add_map_x_26_sg_up), .sg_down(_add_map_x_26_sg_down), .sg_left(_add_map_x_26_sg_left), .sg_right(_add_map_x_26_sg_right), .wall_t_in(_add_map_x_26_wall_t_in), .moto(_add_map_x_26_moto), .up(_add_map_x_26_up), .right(_add_map_x_26_right), .down(_add_map_x_26_down), .left(_add_map_x_26_left), .start(_add_map_x_26_start), .goal(_add_map_x_26_goal), .now(_add_map_x_26_now), .distance(_add_map_x_26_distance));
add_map add_map_x_25 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_25_add_exe), .end_wall(_add_map_x_25_end_wall), .all_s_g(_add_map_x_25_all_s_g), .all_s_g_near(_add_map_x_25_all_s_g_near), .data_out(_add_map_x_25_data_out), .data_out_index(_add_map_x_25_data_out_index), .data_near(_add_map_x_25_data_near), .wall_t_out(_add_map_x_25_wall_t_out), .data_org(_add_map_x_25_data_org), .data_org_near(_add_map_x_25_data_org_near), .s_g(_add_map_x_25_s_g), .s_g_near(_add_map_x_25_s_g_near), .wall_end_in(_add_map_x_25_wall_end_in), .all_sg_up(_add_map_x_25_all_sg_up), .all_sg_down(_add_map_x_25_all_sg_down), .all_sg_right(_add_map_x_25_all_sg_right), .all_sg_left(_add_map_x_25_all_sg_left), .moto_org_near(_add_map_x_25_moto_org_near), .moto_org_near1(_add_map_x_25_moto_org_near1), .moto_org_near2(_add_map_x_25_moto_org_near2), .moto_org_near3(_add_map_x_25_moto_org_near3), .moto_org(_add_map_x_25_moto_org), .sg_up(_add_map_x_25_sg_up), .sg_down(_add_map_x_25_sg_down), .sg_left(_add_map_x_25_sg_left), .sg_right(_add_map_x_25_sg_right), .wall_t_in(_add_map_x_25_wall_t_in), .moto(_add_map_x_25_moto), .up(_add_map_x_25_up), .right(_add_map_x_25_right), .down(_add_map_x_25_down), .left(_add_map_x_25_left), .start(_add_map_x_25_start), .goal(_add_map_x_25_goal), .now(_add_map_x_25_now), .distance(_add_map_x_25_distance));
add_map add_map_x_24 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_24_add_exe), .end_wall(_add_map_x_24_end_wall), .all_s_g(_add_map_x_24_all_s_g), .all_s_g_near(_add_map_x_24_all_s_g_near), .data_out(_add_map_x_24_data_out), .data_out_index(_add_map_x_24_data_out_index), .data_near(_add_map_x_24_data_near), .wall_t_out(_add_map_x_24_wall_t_out), .data_org(_add_map_x_24_data_org), .data_org_near(_add_map_x_24_data_org_near), .s_g(_add_map_x_24_s_g), .s_g_near(_add_map_x_24_s_g_near), .wall_end_in(_add_map_x_24_wall_end_in), .all_sg_up(_add_map_x_24_all_sg_up), .all_sg_down(_add_map_x_24_all_sg_down), .all_sg_right(_add_map_x_24_all_sg_right), .all_sg_left(_add_map_x_24_all_sg_left), .moto_org_near(_add_map_x_24_moto_org_near), .moto_org_near1(_add_map_x_24_moto_org_near1), .moto_org_near2(_add_map_x_24_moto_org_near2), .moto_org_near3(_add_map_x_24_moto_org_near3), .moto_org(_add_map_x_24_moto_org), .sg_up(_add_map_x_24_sg_up), .sg_down(_add_map_x_24_sg_down), .sg_left(_add_map_x_24_sg_left), .sg_right(_add_map_x_24_sg_right), .wall_t_in(_add_map_x_24_wall_t_in), .moto(_add_map_x_24_moto), .up(_add_map_x_24_up), .right(_add_map_x_24_right), .down(_add_map_x_24_down), .left(_add_map_x_24_left), .start(_add_map_x_24_start), .goal(_add_map_x_24_goal), .now(_add_map_x_24_now), .distance(_add_map_x_24_distance));
add_map add_map_x_23 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_23_add_exe), .end_wall(_add_map_x_23_end_wall), .all_s_g(_add_map_x_23_all_s_g), .all_s_g_near(_add_map_x_23_all_s_g_near), .data_out(_add_map_x_23_data_out), .data_out_index(_add_map_x_23_data_out_index), .data_near(_add_map_x_23_data_near), .wall_t_out(_add_map_x_23_wall_t_out), .data_org(_add_map_x_23_data_org), .data_org_near(_add_map_x_23_data_org_near), .s_g(_add_map_x_23_s_g), .s_g_near(_add_map_x_23_s_g_near), .wall_end_in(_add_map_x_23_wall_end_in), .all_sg_up(_add_map_x_23_all_sg_up), .all_sg_down(_add_map_x_23_all_sg_down), .all_sg_right(_add_map_x_23_all_sg_right), .all_sg_left(_add_map_x_23_all_sg_left), .moto_org_near(_add_map_x_23_moto_org_near), .moto_org_near1(_add_map_x_23_moto_org_near1), .moto_org_near2(_add_map_x_23_moto_org_near2), .moto_org_near3(_add_map_x_23_moto_org_near3), .moto_org(_add_map_x_23_moto_org), .sg_up(_add_map_x_23_sg_up), .sg_down(_add_map_x_23_sg_down), .sg_left(_add_map_x_23_sg_left), .sg_right(_add_map_x_23_sg_right), .wall_t_in(_add_map_x_23_wall_t_in), .moto(_add_map_x_23_moto), .up(_add_map_x_23_up), .right(_add_map_x_23_right), .down(_add_map_x_23_down), .left(_add_map_x_23_left), .start(_add_map_x_23_start), .goal(_add_map_x_23_goal), .now(_add_map_x_23_now), .distance(_add_map_x_23_distance));
add_map add_map_x_22 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_22_add_exe), .end_wall(_add_map_x_22_end_wall), .all_s_g(_add_map_x_22_all_s_g), .all_s_g_near(_add_map_x_22_all_s_g_near), .data_out(_add_map_x_22_data_out), .data_out_index(_add_map_x_22_data_out_index), .data_near(_add_map_x_22_data_near), .wall_t_out(_add_map_x_22_wall_t_out), .data_org(_add_map_x_22_data_org), .data_org_near(_add_map_x_22_data_org_near), .s_g(_add_map_x_22_s_g), .s_g_near(_add_map_x_22_s_g_near), .wall_end_in(_add_map_x_22_wall_end_in), .all_sg_up(_add_map_x_22_all_sg_up), .all_sg_down(_add_map_x_22_all_sg_down), .all_sg_right(_add_map_x_22_all_sg_right), .all_sg_left(_add_map_x_22_all_sg_left), .moto_org_near(_add_map_x_22_moto_org_near), .moto_org_near1(_add_map_x_22_moto_org_near1), .moto_org_near2(_add_map_x_22_moto_org_near2), .moto_org_near3(_add_map_x_22_moto_org_near3), .moto_org(_add_map_x_22_moto_org), .sg_up(_add_map_x_22_sg_up), .sg_down(_add_map_x_22_sg_down), .sg_left(_add_map_x_22_sg_left), .sg_right(_add_map_x_22_sg_right), .wall_t_in(_add_map_x_22_wall_t_in), .moto(_add_map_x_22_moto), .up(_add_map_x_22_up), .right(_add_map_x_22_right), .down(_add_map_x_22_down), .left(_add_map_x_22_left), .start(_add_map_x_22_start), .goal(_add_map_x_22_goal), .now(_add_map_x_22_now), .distance(_add_map_x_22_distance));
add_map add_map_x_21 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_21_add_exe), .end_wall(_add_map_x_21_end_wall), .all_s_g(_add_map_x_21_all_s_g), .all_s_g_near(_add_map_x_21_all_s_g_near), .data_out(_add_map_x_21_data_out), .data_out_index(_add_map_x_21_data_out_index), .data_near(_add_map_x_21_data_near), .wall_t_out(_add_map_x_21_wall_t_out), .data_org(_add_map_x_21_data_org), .data_org_near(_add_map_x_21_data_org_near), .s_g(_add_map_x_21_s_g), .s_g_near(_add_map_x_21_s_g_near), .wall_end_in(_add_map_x_21_wall_end_in), .all_sg_up(_add_map_x_21_all_sg_up), .all_sg_down(_add_map_x_21_all_sg_down), .all_sg_right(_add_map_x_21_all_sg_right), .all_sg_left(_add_map_x_21_all_sg_left), .moto_org_near(_add_map_x_21_moto_org_near), .moto_org_near1(_add_map_x_21_moto_org_near1), .moto_org_near2(_add_map_x_21_moto_org_near2), .moto_org_near3(_add_map_x_21_moto_org_near3), .moto_org(_add_map_x_21_moto_org), .sg_up(_add_map_x_21_sg_up), .sg_down(_add_map_x_21_sg_down), .sg_left(_add_map_x_21_sg_left), .sg_right(_add_map_x_21_sg_right), .wall_t_in(_add_map_x_21_wall_t_in), .moto(_add_map_x_21_moto), .up(_add_map_x_21_up), .right(_add_map_x_21_right), .down(_add_map_x_21_down), .left(_add_map_x_21_left), .start(_add_map_x_21_start), .goal(_add_map_x_21_goal), .now(_add_map_x_21_now), .distance(_add_map_x_21_distance));
add_map add_map_x_20 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_20_add_exe), .end_wall(_add_map_x_20_end_wall), .all_s_g(_add_map_x_20_all_s_g), .all_s_g_near(_add_map_x_20_all_s_g_near), .data_out(_add_map_x_20_data_out), .data_out_index(_add_map_x_20_data_out_index), .data_near(_add_map_x_20_data_near), .wall_t_out(_add_map_x_20_wall_t_out), .data_org(_add_map_x_20_data_org), .data_org_near(_add_map_x_20_data_org_near), .s_g(_add_map_x_20_s_g), .s_g_near(_add_map_x_20_s_g_near), .wall_end_in(_add_map_x_20_wall_end_in), .all_sg_up(_add_map_x_20_all_sg_up), .all_sg_down(_add_map_x_20_all_sg_down), .all_sg_right(_add_map_x_20_all_sg_right), .all_sg_left(_add_map_x_20_all_sg_left), .moto_org_near(_add_map_x_20_moto_org_near), .moto_org_near1(_add_map_x_20_moto_org_near1), .moto_org_near2(_add_map_x_20_moto_org_near2), .moto_org_near3(_add_map_x_20_moto_org_near3), .moto_org(_add_map_x_20_moto_org), .sg_up(_add_map_x_20_sg_up), .sg_down(_add_map_x_20_sg_down), .sg_left(_add_map_x_20_sg_left), .sg_right(_add_map_x_20_sg_right), .wall_t_in(_add_map_x_20_wall_t_in), .moto(_add_map_x_20_moto), .up(_add_map_x_20_up), .right(_add_map_x_20_right), .down(_add_map_x_20_down), .left(_add_map_x_20_left), .start(_add_map_x_20_start), .goal(_add_map_x_20_goal), .now(_add_map_x_20_now), .distance(_add_map_x_20_distance));
add_map add_map_x_19 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_19_add_exe), .end_wall(_add_map_x_19_end_wall), .all_s_g(_add_map_x_19_all_s_g), .all_s_g_near(_add_map_x_19_all_s_g_near), .data_out(_add_map_x_19_data_out), .data_out_index(_add_map_x_19_data_out_index), .data_near(_add_map_x_19_data_near), .wall_t_out(_add_map_x_19_wall_t_out), .data_org(_add_map_x_19_data_org), .data_org_near(_add_map_x_19_data_org_near), .s_g(_add_map_x_19_s_g), .s_g_near(_add_map_x_19_s_g_near), .wall_end_in(_add_map_x_19_wall_end_in), .all_sg_up(_add_map_x_19_all_sg_up), .all_sg_down(_add_map_x_19_all_sg_down), .all_sg_right(_add_map_x_19_all_sg_right), .all_sg_left(_add_map_x_19_all_sg_left), .moto_org_near(_add_map_x_19_moto_org_near), .moto_org_near1(_add_map_x_19_moto_org_near1), .moto_org_near2(_add_map_x_19_moto_org_near2), .moto_org_near3(_add_map_x_19_moto_org_near3), .moto_org(_add_map_x_19_moto_org), .sg_up(_add_map_x_19_sg_up), .sg_down(_add_map_x_19_sg_down), .sg_left(_add_map_x_19_sg_left), .sg_right(_add_map_x_19_sg_right), .wall_t_in(_add_map_x_19_wall_t_in), .moto(_add_map_x_19_moto), .up(_add_map_x_19_up), .right(_add_map_x_19_right), .down(_add_map_x_19_down), .left(_add_map_x_19_left), .start(_add_map_x_19_start), .goal(_add_map_x_19_goal), .now(_add_map_x_19_now), .distance(_add_map_x_19_distance));
add_map add_map_x_18 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_18_add_exe), .end_wall(_add_map_x_18_end_wall), .all_s_g(_add_map_x_18_all_s_g), .all_s_g_near(_add_map_x_18_all_s_g_near), .data_out(_add_map_x_18_data_out), .data_out_index(_add_map_x_18_data_out_index), .data_near(_add_map_x_18_data_near), .wall_t_out(_add_map_x_18_wall_t_out), .data_org(_add_map_x_18_data_org), .data_org_near(_add_map_x_18_data_org_near), .s_g(_add_map_x_18_s_g), .s_g_near(_add_map_x_18_s_g_near), .wall_end_in(_add_map_x_18_wall_end_in), .all_sg_up(_add_map_x_18_all_sg_up), .all_sg_down(_add_map_x_18_all_sg_down), .all_sg_right(_add_map_x_18_all_sg_right), .all_sg_left(_add_map_x_18_all_sg_left), .moto_org_near(_add_map_x_18_moto_org_near), .moto_org_near1(_add_map_x_18_moto_org_near1), .moto_org_near2(_add_map_x_18_moto_org_near2), .moto_org_near3(_add_map_x_18_moto_org_near3), .moto_org(_add_map_x_18_moto_org), .sg_up(_add_map_x_18_sg_up), .sg_down(_add_map_x_18_sg_down), .sg_left(_add_map_x_18_sg_left), .sg_right(_add_map_x_18_sg_right), .wall_t_in(_add_map_x_18_wall_t_in), .moto(_add_map_x_18_moto), .up(_add_map_x_18_up), .right(_add_map_x_18_right), .down(_add_map_x_18_down), .left(_add_map_x_18_left), .start(_add_map_x_18_start), .goal(_add_map_x_18_goal), .now(_add_map_x_18_now), .distance(_add_map_x_18_distance));
add_map add_map_x_17 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_17_add_exe), .end_wall(_add_map_x_17_end_wall), .all_s_g(_add_map_x_17_all_s_g), .all_s_g_near(_add_map_x_17_all_s_g_near), .data_out(_add_map_x_17_data_out), .data_out_index(_add_map_x_17_data_out_index), .data_near(_add_map_x_17_data_near), .wall_t_out(_add_map_x_17_wall_t_out), .data_org(_add_map_x_17_data_org), .data_org_near(_add_map_x_17_data_org_near), .s_g(_add_map_x_17_s_g), .s_g_near(_add_map_x_17_s_g_near), .wall_end_in(_add_map_x_17_wall_end_in), .all_sg_up(_add_map_x_17_all_sg_up), .all_sg_down(_add_map_x_17_all_sg_down), .all_sg_right(_add_map_x_17_all_sg_right), .all_sg_left(_add_map_x_17_all_sg_left), .moto_org_near(_add_map_x_17_moto_org_near), .moto_org_near1(_add_map_x_17_moto_org_near1), .moto_org_near2(_add_map_x_17_moto_org_near2), .moto_org_near3(_add_map_x_17_moto_org_near3), .moto_org(_add_map_x_17_moto_org), .sg_up(_add_map_x_17_sg_up), .sg_down(_add_map_x_17_sg_down), .sg_left(_add_map_x_17_sg_left), .sg_right(_add_map_x_17_sg_right), .wall_t_in(_add_map_x_17_wall_t_in), .moto(_add_map_x_17_moto), .up(_add_map_x_17_up), .right(_add_map_x_17_right), .down(_add_map_x_17_down), .left(_add_map_x_17_left), .start(_add_map_x_17_start), .goal(_add_map_x_17_goal), .now(_add_map_x_17_now), .distance(_add_map_x_17_distance));
add_map add_map_x_16 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_16_add_exe), .end_wall(_add_map_x_16_end_wall), .all_s_g(_add_map_x_16_all_s_g), .all_s_g_near(_add_map_x_16_all_s_g_near), .data_out(_add_map_x_16_data_out), .data_out_index(_add_map_x_16_data_out_index), .data_near(_add_map_x_16_data_near), .wall_t_out(_add_map_x_16_wall_t_out), .data_org(_add_map_x_16_data_org), .data_org_near(_add_map_x_16_data_org_near), .s_g(_add_map_x_16_s_g), .s_g_near(_add_map_x_16_s_g_near), .wall_end_in(_add_map_x_16_wall_end_in), .all_sg_up(_add_map_x_16_all_sg_up), .all_sg_down(_add_map_x_16_all_sg_down), .all_sg_right(_add_map_x_16_all_sg_right), .all_sg_left(_add_map_x_16_all_sg_left), .moto_org_near(_add_map_x_16_moto_org_near), .moto_org_near1(_add_map_x_16_moto_org_near1), .moto_org_near2(_add_map_x_16_moto_org_near2), .moto_org_near3(_add_map_x_16_moto_org_near3), .moto_org(_add_map_x_16_moto_org), .sg_up(_add_map_x_16_sg_up), .sg_down(_add_map_x_16_sg_down), .sg_left(_add_map_x_16_sg_left), .sg_right(_add_map_x_16_sg_right), .wall_t_in(_add_map_x_16_wall_t_in), .moto(_add_map_x_16_moto), .up(_add_map_x_16_up), .right(_add_map_x_16_right), .down(_add_map_x_16_down), .left(_add_map_x_16_left), .start(_add_map_x_16_start), .goal(_add_map_x_16_goal), .now(_add_map_x_16_now), .distance(_add_map_x_16_distance));
add_map add_map_x_15 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_15_add_exe), .end_wall(_add_map_x_15_end_wall), .all_s_g(_add_map_x_15_all_s_g), .all_s_g_near(_add_map_x_15_all_s_g_near), .data_out(_add_map_x_15_data_out), .data_out_index(_add_map_x_15_data_out_index), .data_near(_add_map_x_15_data_near), .wall_t_out(_add_map_x_15_wall_t_out), .data_org(_add_map_x_15_data_org), .data_org_near(_add_map_x_15_data_org_near), .s_g(_add_map_x_15_s_g), .s_g_near(_add_map_x_15_s_g_near), .wall_end_in(_add_map_x_15_wall_end_in), .all_sg_up(_add_map_x_15_all_sg_up), .all_sg_down(_add_map_x_15_all_sg_down), .all_sg_right(_add_map_x_15_all_sg_right), .all_sg_left(_add_map_x_15_all_sg_left), .moto_org_near(_add_map_x_15_moto_org_near), .moto_org_near1(_add_map_x_15_moto_org_near1), .moto_org_near2(_add_map_x_15_moto_org_near2), .moto_org_near3(_add_map_x_15_moto_org_near3), .moto_org(_add_map_x_15_moto_org), .sg_up(_add_map_x_15_sg_up), .sg_down(_add_map_x_15_sg_down), .sg_left(_add_map_x_15_sg_left), .sg_right(_add_map_x_15_sg_right), .wall_t_in(_add_map_x_15_wall_t_in), .moto(_add_map_x_15_moto), .up(_add_map_x_15_up), .right(_add_map_x_15_right), .down(_add_map_x_15_down), .left(_add_map_x_15_left), .start(_add_map_x_15_start), .goal(_add_map_x_15_goal), .now(_add_map_x_15_now), .distance(_add_map_x_15_distance));
add_map add_map_x_14 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_14_add_exe), .end_wall(_add_map_x_14_end_wall), .all_s_g(_add_map_x_14_all_s_g), .all_s_g_near(_add_map_x_14_all_s_g_near), .data_out(_add_map_x_14_data_out), .data_out_index(_add_map_x_14_data_out_index), .data_near(_add_map_x_14_data_near), .wall_t_out(_add_map_x_14_wall_t_out), .data_org(_add_map_x_14_data_org), .data_org_near(_add_map_x_14_data_org_near), .s_g(_add_map_x_14_s_g), .s_g_near(_add_map_x_14_s_g_near), .wall_end_in(_add_map_x_14_wall_end_in), .all_sg_up(_add_map_x_14_all_sg_up), .all_sg_down(_add_map_x_14_all_sg_down), .all_sg_right(_add_map_x_14_all_sg_right), .all_sg_left(_add_map_x_14_all_sg_left), .moto_org_near(_add_map_x_14_moto_org_near), .moto_org_near1(_add_map_x_14_moto_org_near1), .moto_org_near2(_add_map_x_14_moto_org_near2), .moto_org_near3(_add_map_x_14_moto_org_near3), .moto_org(_add_map_x_14_moto_org), .sg_up(_add_map_x_14_sg_up), .sg_down(_add_map_x_14_sg_down), .sg_left(_add_map_x_14_sg_left), .sg_right(_add_map_x_14_sg_right), .wall_t_in(_add_map_x_14_wall_t_in), .moto(_add_map_x_14_moto), .up(_add_map_x_14_up), .right(_add_map_x_14_right), .down(_add_map_x_14_down), .left(_add_map_x_14_left), .start(_add_map_x_14_start), .goal(_add_map_x_14_goal), .now(_add_map_x_14_now), .distance(_add_map_x_14_distance));
add_map add_map_x_13 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_13_add_exe), .end_wall(_add_map_x_13_end_wall), .all_s_g(_add_map_x_13_all_s_g), .all_s_g_near(_add_map_x_13_all_s_g_near), .data_out(_add_map_x_13_data_out), .data_out_index(_add_map_x_13_data_out_index), .data_near(_add_map_x_13_data_near), .wall_t_out(_add_map_x_13_wall_t_out), .data_org(_add_map_x_13_data_org), .data_org_near(_add_map_x_13_data_org_near), .s_g(_add_map_x_13_s_g), .s_g_near(_add_map_x_13_s_g_near), .wall_end_in(_add_map_x_13_wall_end_in), .all_sg_up(_add_map_x_13_all_sg_up), .all_sg_down(_add_map_x_13_all_sg_down), .all_sg_right(_add_map_x_13_all_sg_right), .all_sg_left(_add_map_x_13_all_sg_left), .moto_org_near(_add_map_x_13_moto_org_near), .moto_org_near1(_add_map_x_13_moto_org_near1), .moto_org_near2(_add_map_x_13_moto_org_near2), .moto_org_near3(_add_map_x_13_moto_org_near3), .moto_org(_add_map_x_13_moto_org), .sg_up(_add_map_x_13_sg_up), .sg_down(_add_map_x_13_sg_down), .sg_left(_add_map_x_13_sg_left), .sg_right(_add_map_x_13_sg_right), .wall_t_in(_add_map_x_13_wall_t_in), .moto(_add_map_x_13_moto), .up(_add_map_x_13_up), .right(_add_map_x_13_right), .down(_add_map_x_13_down), .left(_add_map_x_13_left), .start(_add_map_x_13_start), .goal(_add_map_x_13_goal), .now(_add_map_x_13_now), .distance(_add_map_x_13_distance));
add_map add_map_x_12 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_12_add_exe), .end_wall(_add_map_x_12_end_wall), .all_s_g(_add_map_x_12_all_s_g), .all_s_g_near(_add_map_x_12_all_s_g_near), .data_out(_add_map_x_12_data_out), .data_out_index(_add_map_x_12_data_out_index), .data_near(_add_map_x_12_data_near), .wall_t_out(_add_map_x_12_wall_t_out), .data_org(_add_map_x_12_data_org), .data_org_near(_add_map_x_12_data_org_near), .s_g(_add_map_x_12_s_g), .s_g_near(_add_map_x_12_s_g_near), .wall_end_in(_add_map_x_12_wall_end_in), .all_sg_up(_add_map_x_12_all_sg_up), .all_sg_down(_add_map_x_12_all_sg_down), .all_sg_right(_add_map_x_12_all_sg_right), .all_sg_left(_add_map_x_12_all_sg_left), .moto_org_near(_add_map_x_12_moto_org_near), .moto_org_near1(_add_map_x_12_moto_org_near1), .moto_org_near2(_add_map_x_12_moto_org_near2), .moto_org_near3(_add_map_x_12_moto_org_near3), .moto_org(_add_map_x_12_moto_org), .sg_up(_add_map_x_12_sg_up), .sg_down(_add_map_x_12_sg_down), .sg_left(_add_map_x_12_sg_left), .sg_right(_add_map_x_12_sg_right), .wall_t_in(_add_map_x_12_wall_t_in), .moto(_add_map_x_12_moto), .up(_add_map_x_12_up), .right(_add_map_x_12_right), .down(_add_map_x_12_down), .left(_add_map_x_12_left), .start(_add_map_x_12_start), .goal(_add_map_x_12_goal), .now(_add_map_x_12_now), .distance(_add_map_x_12_distance));
add_map add_map_x_11 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_11_add_exe), .end_wall(_add_map_x_11_end_wall), .all_s_g(_add_map_x_11_all_s_g), .all_s_g_near(_add_map_x_11_all_s_g_near), .data_out(_add_map_x_11_data_out), .data_out_index(_add_map_x_11_data_out_index), .data_near(_add_map_x_11_data_near), .wall_t_out(_add_map_x_11_wall_t_out), .data_org(_add_map_x_11_data_org), .data_org_near(_add_map_x_11_data_org_near), .s_g(_add_map_x_11_s_g), .s_g_near(_add_map_x_11_s_g_near), .wall_end_in(_add_map_x_11_wall_end_in), .all_sg_up(_add_map_x_11_all_sg_up), .all_sg_down(_add_map_x_11_all_sg_down), .all_sg_right(_add_map_x_11_all_sg_right), .all_sg_left(_add_map_x_11_all_sg_left), .moto_org_near(_add_map_x_11_moto_org_near), .moto_org_near1(_add_map_x_11_moto_org_near1), .moto_org_near2(_add_map_x_11_moto_org_near2), .moto_org_near3(_add_map_x_11_moto_org_near3), .moto_org(_add_map_x_11_moto_org), .sg_up(_add_map_x_11_sg_up), .sg_down(_add_map_x_11_sg_down), .sg_left(_add_map_x_11_sg_left), .sg_right(_add_map_x_11_sg_right), .wall_t_in(_add_map_x_11_wall_t_in), .moto(_add_map_x_11_moto), .up(_add_map_x_11_up), .right(_add_map_x_11_right), .down(_add_map_x_11_down), .left(_add_map_x_11_left), .start(_add_map_x_11_start), .goal(_add_map_x_11_goal), .now(_add_map_x_11_now), .distance(_add_map_x_11_distance));
add_map add_map_x_10 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_10_add_exe), .end_wall(_add_map_x_10_end_wall), .all_s_g(_add_map_x_10_all_s_g), .all_s_g_near(_add_map_x_10_all_s_g_near), .data_out(_add_map_x_10_data_out), .data_out_index(_add_map_x_10_data_out_index), .data_near(_add_map_x_10_data_near), .wall_t_out(_add_map_x_10_wall_t_out), .data_org(_add_map_x_10_data_org), .data_org_near(_add_map_x_10_data_org_near), .s_g(_add_map_x_10_s_g), .s_g_near(_add_map_x_10_s_g_near), .wall_end_in(_add_map_x_10_wall_end_in), .all_sg_up(_add_map_x_10_all_sg_up), .all_sg_down(_add_map_x_10_all_sg_down), .all_sg_right(_add_map_x_10_all_sg_right), .all_sg_left(_add_map_x_10_all_sg_left), .moto_org_near(_add_map_x_10_moto_org_near), .moto_org_near1(_add_map_x_10_moto_org_near1), .moto_org_near2(_add_map_x_10_moto_org_near2), .moto_org_near3(_add_map_x_10_moto_org_near3), .moto_org(_add_map_x_10_moto_org), .sg_up(_add_map_x_10_sg_up), .sg_down(_add_map_x_10_sg_down), .sg_left(_add_map_x_10_sg_left), .sg_right(_add_map_x_10_sg_right), .wall_t_in(_add_map_x_10_wall_t_in), .moto(_add_map_x_10_moto), .up(_add_map_x_10_up), .right(_add_map_x_10_right), .down(_add_map_x_10_down), .left(_add_map_x_10_left), .start(_add_map_x_10_start), .goal(_add_map_x_10_goal), .now(_add_map_x_10_now), .distance(_add_map_x_10_distance));
add_map add_map_x_9 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_9_add_exe), .end_wall(_add_map_x_9_end_wall), .all_s_g(_add_map_x_9_all_s_g), .all_s_g_near(_add_map_x_9_all_s_g_near), .data_out(_add_map_x_9_data_out), .data_out_index(_add_map_x_9_data_out_index), .data_near(_add_map_x_9_data_near), .wall_t_out(_add_map_x_9_wall_t_out), .data_org(_add_map_x_9_data_org), .data_org_near(_add_map_x_9_data_org_near), .s_g(_add_map_x_9_s_g), .s_g_near(_add_map_x_9_s_g_near), .wall_end_in(_add_map_x_9_wall_end_in), .all_sg_up(_add_map_x_9_all_sg_up), .all_sg_down(_add_map_x_9_all_sg_down), .all_sg_right(_add_map_x_9_all_sg_right), .all_sg_left(_add_map_x_9_all_sg_left), .moto_org_near(_add_map_x_9_moto_org_near), .moto_org_near1(_add_map_x_9_moto_org_near1), .moto_org_near2(_add_map_x_9_moto_org_near2), .moto_org_near3(_add_map_x_9_moto_org_near3), .moto_org(_add_map_x_9_moto_org), .sg_up(_add_map_x_9_sg_up), .sg_down(_add_map_x_9_sg_down), .sg_left(_add_map_x_9_sg_left), .sg_right(_add_map_x_9_sg_right), .wall_t_in(_add_map_x_9_wall_t_in), .moto(_add_map_x_9_moto), .up(_add_map_x_9_up), .right(_add_map_x_9_right), .down(_add_map_x_9_down), .left(_add_map_x_9_left), .start(_add_map_x_9_start), .goal(_add_map_x_9_goal), .now(_add_map_x_9_now), .distance(_add_map_x_9_distance));
add_map add_map_x_8 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_8_add_exe), .end_wall(_add_map_x_8_end_wall), .all_s_g(_add_map_x_8_all_s_g), .all_s_g_near(_add_map_x_8_all_s_g_near), .data_out(_add_map_x_8_data_out), .data_out_index(_add_map_x_8_data_out_index), .data_near(_add_map_x_8_data_near), .wall_t_out(_add_map_x_8_wall_t_out), .data_org(_add_map_x_8_data_org), .data_org_near(_add_map_x_8_data_org_near), .s_g(_add_map_x_8_s_g), .s_g_near(_add_map_x_8_s_g_near), .wall_end_in(_add_map_x_8_wall_end_in), .all_sg_up(_add_map_x_8_all_sg_up), .all_sg_down(_add_map_x_8_all_sg_down), .all_sg_right(_add_map_x_8_all_sg_right), .all_sg_left(_add_map_x_8_all_sg_left), .moto_org_near(_add_map_x_8_moto_org_near), .moto_org_near1(_add_map_x_8_moto_org_near1), .moto_org_near2(_add_map_x_8_moto_org_near2), .moto_org_near3(_add_map_x_8_moto_org_near3), .moto_org(_add_map_x_8_moto_org), .sg_up(_add_map_x_8_sg_up), .sg_down(_add_map_x_8_sg_down), .sg_left(_add_map_x_8_sg_left), .sg_right(_add_map_x_8_sg_right), .wall_t_in(_add_map_x_8_wall_t_in), .moto(_add_map_x_8_moto), .up(_add_map_x_8_up), .right(_add_map_x_8_right), .down(_add_map_x_8_down), .left(_add_map_x_8_left), .start(_add_map_x_8_start), .goal(_add_map_x_8_goal), .now(_add_map_x_8_now), .distance(_add_map_x_8_distance));
add_map add_map_x_7 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_7_add_exe), .end_wall(_add_map_x_7_end_wall), .all_s_g(_add_map_x_7_all_s_g), .all_s_g_near(_add_map_x_7_all_s_g_near), .data_out(_add_map_x_7_data_out), .data_out_index(_add_map_x_7_data_out_index), .data_near(_add_map_x_7_data_near), .wall_t_out(_add_map_x_7_wall_t_out), .data_org(_add_map_x_7_data_org), .data_org_near(_add_map_x_7_data_org_near), .s_g(_add_map_x_7_s_g), .s_g_near(_add_map_x_7_s_g_near), .wall_end_in(_add_map_x_7_wall_end_in), .all_sg_up(_add_map_x_7_all_sg_up), .all_sg_down(_add_map_x_7_all_sg_down), .all_sg_right(_add_map_x_7_all_sg_right), .all_sg_left(_add_map_x_7_all_sg_left), .moto_org_near(_add_map_x_7_moto_org_near), .moto_org_near1(_add_map_x_7_moto_org_near1), .moto_org_near2(_add_map_x_7_moto_org_near2), .moto_org_near3(_add_map_x_7_moto_org_near3), .moto_org(_add_map_x_7_moto_org), .sg_up(_add_map_x_7_sg_up), .sg_down(_add_map_x_7_sg_down), .sg_left(_add_map_x_7_sg_left), .sg_right(_add_map_x_7_sg_right), .wall_t_in(_add_map_x_7_wall_t_in), .moto(_add_map_x_7_moto), .up(_add_map_x_7_up), .right(_add_map_x_7_right), .down(_add_map_x_7_down), .left(_add_map_x_7_left), .start(_add_map_x_7_start), .goal(_add_map_x_7_goal), .now(_add_map_x_7_now), .distance(_add_map_x_7_distance));
add_map add_map_x_6 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_6_add_exe), .end_wall(_add_map_x_6_end_wall), .all_s_g(_add_map_x_6_all_s_g), .all_s_g_near(_add_map_x_6_all_s_g_near), .data_out(_add_map_x_6_data_out), .data_out_index(_add_map_x_6_data_out_index), .data_near(_add_map_x_6_data_near), .wall_t_out(_add_map_x_6_wall_t_out), .data_org(_add_map_x_6_data_org), .data_org_near(_add_map_x_6_data_org_near), .s_g(_add_map_x_6_s_g), .s_g_near(_add_map_x_6_s_g_near), .wall_end_in(_add_map_x_6_wall_end_in), .all_sg_up(_add_map_x_6_all_sg_up), .all_sg_down(_add_map_x_6_all_sg_down), .all_sg_right(_add_map_x_6_all_sg_right), .all_sg_left(_add_map_x_6_all_sg_left), .moto_org_near(_add_map_x_6_moto_org_near), .moto_org_near1(_add_map_x_6_moto_org_near1), .moto_org_near2(_add_map_x_6_moto_org_near2), .moto_org_near3(_add_map_x_6_moto_org_near3), .moto_org(_add_map_x_6_moto_org), .sg_up(_add_map_x_6_sg_up), .sg_down(_add_map_x_6_sg_down), .sg_left(_add_map_x_6_sg_left), .sg_right(_add_map_x_6_sg_right), .wall_t_in(_add_map_x_6_wall_t_in), .moto(_add_map_x_6_moto), .up(_add_map_x_6_up), .right(_add_map_x_6_right), .down(_add_map_x_6_down), .left(_add_map_x_6_left), .start(_add_map_x_6_start), .goal(_add_map_x_6_goal), .now(_add_map_x_6_now), .distance(_add_map_x_6_distance));
add_map add_map_x_5 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_5_add_exe), .end_wall(_add_map_x_5_end_wall), .all_s_g(_add_map_x_5_all_s_g), .all_s_g_near(_add_map_x_5_all_s_g_near), .data_out(_add_map_x_5_data_out), .data_out_index(_add_map_x_5_data_out_index), .data_near(_add_map_x_5_data_near), .wall_t_out(_add_map_x_5_wall_t_out), .data_org(_add_map_x_5_data_org), .data_org_near(_add_map_x_5_data_org_near), .s_g(_add_map_x_5_s_g), .s_g_near(_add_map_x_5_s_g_near), .wall_end_in(_add_map_x_5_wall_end_in), .all_sg_up(_add_map_x_5_all_sg_up), .all_sg_down(_add_map_x_5_all_sg_down), .all_sg_right(_add_map_x_5_all_sg_right), .all_sg_left(_add_map_x_5_all_sg_left), .moto_org_near(_add_map_x_5_moto_org_near), .moto_org_near1(_add_map_x_5_moto_org_near1), .moto_org_near2(_add_map_x_5_moto_org_near2), .moto_org_near3(_add_map_x_5_moto_org_near3), .moto_org(_add_map_x_5_moto_org), .sg_up(_add_map_x_5_sg_up), .sg_down(_add_map_x_5_sg_down), .sg_left(_add_map_x_5_sg_left), .sg_right(_add_map_x_5_sg_right), .wall_t_in(_add_map_x_5_wall_t_in), .moto(_add_map_x_5_moto), .up(_add_map_x_5_up), .right(_add_map_x_5_right), .down(_add_map_x_5_down), .left(_add_map_x_5_left), .start(_add_map_x_5_start), .goal(_add_map_x_5_goal), .now(_add_map_x_5_now), .distance(_add_map_x_5_distance));
add_map add_map_x_4 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_4_add_exe), .end_wall(_add_map_x_4_end_wall), .all_s_g(_add_map_x_4_all_s_g), .all_s_g_near(_add_map_x_4_all_s_g_near), .data_out(_add_map_x_4_data_out), .data_out_index(_add_map_x_4_data_out_index), .data_near(_add_map_x_4_data_near), .wall_t_out(_add_map_x_4_wall_t_out), .data_org(_add_map_x_4_data_org), .data_org_near(_add_map_x_4_data_org_near), .s_g(_add_map_x_4_s_g), .s_g_near(_add_map_x_4_s_g_near), .wall_end_in(_add_map_x_4_wall_end_in), .all_sg_up(_add_map_x_4_all_sg_up), .all_sg_down(_add_map_x_4_all_sg_down), .all_sg_right(_add_map_x_4_all_sg_right), .all_sg_left(_add_map_x_4_all_sg_left), .moto_org_near(_add_map_x_4_moto_org_near), .moto_org_near1(_add_map_x_4_moto_org_near1), .moto_org_near2(_add_map_x_4_moto_org_near2), .moto_org_near3(_add_map_x_4_moto_org_near3), .moto_org(_add_map_x_4_moto_org), .sg_up(_add_map_x_4_sg_up), .sg_down(_add_map_x_4_sg_down), .sg_left(_add_map_x_4_sg_left), .sg_right(_add_map_x_4_sg_right), .wall_t_in(_add_map_x_4_wall_t_in), .moto(_add_map_x_4_moto), .up(_add_map_x_4_up), .right(_add_map_x_4_right), .down(_add_map_x_4_down), .left(_add_map_x_4_left), .start(_add_map_x_4_start), .goal(_add_map_x_4_goal), .now(_add_map_x_4_now), .distance(_add_map_x_4_distance));
add_map add_map_x_3 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_3_add_exe), .end_wall(_add_map_x_3_end_wall), .all_s_g(_add_map_x_3_all_s_g), .all_s_g_near(_add_map_x_3_all_s_g_near), .data_out(_add_map_x_3_data_out), .data_out_index(_add_map_x_3_data_out_index), .data_near(_add_map_x_3_data_near), .wall_t_out(_add_map_x_3_wall_t_out), .data_org(_add_map_x_3_data_org), .data_org_near(_add_map_x_3_data_org_near), .s_g(_add_map_x_3_s_g), .s_g_near(_add_map_x_3_s_g_near), .wall_end_in(_add_map_x_3_wall_end_in), .all_sg_up(_add_map_x_3_all_sg_up), .all_sg_down(_add_map_x_3_all_sg_down), .all_sg_right(_add_map_x_3_all_sg_right), .all_sg_left(_add_map_x_3_all_sg_left), .moto_org_near(_add_map_x_3_moto_org_near), .moto_org_near1(_add_map_x_3_moto_org_near1), .moto_org_near2(_add_map_x_3_moto_org_near2), .moto_org_near3(_add_map_x_3_moto_org_near3), .moto_org(_add_map_x_3_moto_org), .sg_up(_add_map_x_3_sg_up), .sg_down(_add_map_x_3_sg_down), .sg_left(_add_map_x_3_sg_left), .sg_right(_add_map_x_3_sg_right), .wall_t_in(_add_map_x_3_wall_t_in), .moto(_add_map_x_3_moto), .up(_add_map_x_3_up), .right(_add_map_x_3_right), .down(_add_map_x_3_down), .left(_add_map_x_3_left), .start(_add_map_x_3_start), .goal(_add_map_x_3_goal), .now(_add_map_x_3_now), .distance(_add_map_x_3_distance));
add_map add_map_x_2 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_2_add_exe), .end_wall(_add_map_x_2_end_wall), .all_s_g(_add_map_x_2_all_s_g), .all_s_g_near(_add_map_x_2_all_s_g_near), .data_out(_add_map_x_2_data_out), .data_out_index(_add_map_x_2_data_out_index), .data_near(_add_map_x_2_data_near), .wall_t_out(_add_map_x_2_wall_t_out), .data_org(_add_map_x_2_data_org), .data_org_near(_add_map_x_2_data_org_near), .s_g(_add_map_x_2_s_g), .s_g_near(_add_map_x_2_s_g_near), .wall_end_in(_add_map_x_2_wall_end_in), .all_sg_up(_add_map_x_2_all_sg_up), .all_sg_down(_add_map_x_2_all_sg_down), .all_sg_right(_add_map_x_2_all_sg_right), .all_sg_left(_add_map_x_2_all_sg_left), .moto_org_near(_add_map_x_2_moto_org_near), .moto_org_near1(_add_map_x_2_moto_org_near1), .moto_org_near2(_add_map_x_2_moto_org_near2), .moto_org_near3(_add_map_x_2_moto_org_near3), .moto_org(_add_map_x_2_moto_org), .sg_up(_add_map_x_2_sg_up), .sg_down(_add_map_x_2_sg_down), .sg_left(_add_map_x_2_sg_left), .sg_right(_add_map_x_2_sg_right), .wall_t_in(_add_map_x_2_wall_t_in), .moto(_add_map_x_2_moto), .up(_add_map_x_2_up), .right(_add_map_x_2_right), .down(_add_map_x_2_down), .left(_add_map_x_2_left), .start(_add_map_x_2_start), .goal(_add_map_x_2_goal), .now(_add_map_x_2_now), .distance(_add_map_x_2_distance));
add_map add_map_x_1 (.m_clock(m_clock), .p_reset( p_reset), .add_exe(_add_map_x_1_add_exe), .end_wall(_add_map_x_1_end_wall), .all_s_g(_add_map_x_1_all_s_g), .all_s_g_near(_add_map_x_1_all_s_g_near), .data_out(_add_map_x_1_data_out), .data_out_index(_add_map_x_1_data_out_index), .data_near(_add_map_x_1_data_near), .wall_t_out(_add_map_x_1_wall_t_out), .data_org(_add_map_x_1_data_org), .data_org_near(_add_map_x_1_data_org_near), .s_g(_add_map_x_1_s_g), .s_g_near(_add_map_x_1_s_g_near), .wall_end_in(_add_map_x_1_wall_end_in), .all_sg_up(_add_map_x_1_all_sg_up), .all_sg_down(_add_map_x_1_all_sg_down), .all_sg_right(_add_map_x_1_all_sg_right), .all_sg_left(_add_map_x_1_all_sg_left), .moto_org_near(_add_map_x_1_moto_org_near), .moto_org_near1(_add_map_x_1_moto_org_near1), .moto_org_near2(_add_map_x_1_moto_org_near2), .moto_org_near3(_add_map_x_1_moto_org_near3), .moto_org(_add_map_x_1_moto_org), .sg_up(_add_map_x_1_sg_up), .sg_down(_add_map_x_1_sg_down), .sg_left(_add_map_x_1_sg_left), .sg_right(_add_map_x_1_sg_right), .wall_t_in(_add_map_x_1_wall_t_in), .moto(_add_map_x_1_moto), .up(_add_map_x_1_up), .right(_add_map_x_1_right), .down(_add_map_x_1_down), .left(_add_map_x_1_left), .start(_add_map_x_1_start), .goal(_add_map_x_1_goal), .now(_add_map_x_1_now), .distance(_add_map_x_1_distance));


// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in33:128'b0)|
    (((in_do&_net_2))?all_sg_in17:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in18:128'b0)|
    (((in_do&_net_2))?all_sg_in19:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)|
    (((in_do&_net_2))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)|
    (((in_do&_net_2))?all_sg_in34:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org18:8'b0)|
    (((in_do&_net_2))?data_in_org17:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?data_in_org19:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org33:8'b0)|
    (((in_do&_net_2))?data_in_org34:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org17:8'b0)|
    (((in_do&_net_2))?data_in_org18:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in18:2'b0)|
    (((in_do&_net_2))?sg_in17:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?2'b00:2'b0)|
    (((in_do&_net_2))?sg_in19:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in33:2'b0)|
    (((in_do&_net_2))?sg_in34:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?2'b00:2'b0)|
    (((in_do&_net_2))?2'b00:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in17:8'b0)|
    (((in_do&_net_2))?data_in18:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in18:8'b0)|
    (((in_do&_net_2))?data_in17:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?data_in19:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in33:8'b0)|
    (((in_do&_net_2))?data_in34:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b00010001:8'b0)|
    (((in_do&_net_2))?8'b00010010:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 97 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 50 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_add_exe)
  begin
#1 if (_add_map_x_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 97 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 50 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_p_reset = p_reset;
   assign  _add_map_x_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in109:128'b0)|
    (((in_do&_net_2))?all_sg_in110:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)|
    (((in_do&_net_2))?all_sg_in108:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in94:128'b0)|
    (((in_do&_net_2))?all_sg_in93:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)|
    (((in_do&_net_2))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org109:8'b0)|
    (((in_do&_net_2))?data_in_org110:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?data_in_org108:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org94:8'b0)|
    (((in_do&_net_2))?data_in_org93:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org110:8'b0)|
    (((in_do&_net_2))?data_in_org109:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in109:2'b0)|
    (((in_do&_net_2))?sg_in110:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?2'b00:2'b0)|
    (((in_do&_net_2))?sg_in108:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?2'b00:2'b0)|
    (((in_do&_net_2))?2'b00:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in94:2'b0)|
    (((in_do&_net_2))?sg_in93:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in110:8'b0)|
    (((in_do&_net_2))?data_in109:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in109:8'b0)|
    (((in_do&_net_2))?data_in110:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?data_in108:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in94:8'b0)|
    (((in_do&_net_2))?data_in93:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b01101110:8'b0)|
    (((in_do&_net_2))?8'b01101101:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_41_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 138 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 91 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_41_add_exe)
  begin
#1 if (_add_map_x_41_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_41_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 138 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 91 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_41_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_41_p_reset = p_reset;
   assign  _add_map_x_41_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in107:128'b0)|
    (((in_do&_net_2))?all_sg_in108:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in109:128'b0)|
    (((in_do&_net_2))?all_sg_in106:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in92:128'b0)|
    (((in_do&_net_2))?all_sg_in91:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)|
    (((in_do&_net_2))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org107:8'b0)|
    (((in_do&_net_2))?data_in_org108:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org109:8'b0)|
    (((in_do&_net_2))?data_in_org106:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org92:8'b0)|
    (((in_do&_net_2))?data_in_org91:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org108:8'b0)|
    (((in_do&_net_2))?data_in_org107:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in107:2'b0)|
    (((in_do&_net_2))?sg_in108:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in109:2'b0)|
    (((in_do&_net_2))?sg_in106:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?2'b00:2'b0)|
    (((in_do&_net_2))?2'b00:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in92:2'b0)|
    (((in_do&_net_2))?sg_in91:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in108:8'b0)|
    (((in_do&_net_2))?data_in107:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in107:8'b0)|
    (((in_do&_net_2))?data_in108:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in109:8'b0)|
    (((in_do&_net_2))?data_in106:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in92:8'b0)|
    (((in_do&_net_2))?data_in91:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b01101100:8'b0)|
    (((in_do&_net_2))?8'b01101011:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_40_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 137 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 90 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_40_add_exe)
  begin
#1 if (_add_map_x_40_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_40_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 137 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 90 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_40_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_40_p_reset = p_reset;
   assign  _add_map_x_40_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in105:128'b0)|
    (((in_do&_net_2))?all_sg_in106:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in107:128'b0)|
    (((in_do&_net_2))?all_sg_in104:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in90:128'b0)|
    (((in_do&_net_2))?all_sg_in89:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)|
    (((in_do&_net_2))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org105:8'b0)|
    (((in_do&_net_2))?data_in_org106:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org107:8'b0)|
    (((in_do&_net_2))?data_in_org104:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org90:8'b0)|
    (((in_do&_net_2))?data_in_org89:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org106:8'b0)|
    (((in_do&_net_2))?data_in_org105:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in105:2'b0)|
    (((in_do&_net_2))?sg_in106:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in107:2'b0)|
    (((in_do&_net_2))?sg_in104:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?2'b00:2'b0)|
    (((in_do&_net_2))?2'b00:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in90:2'b0)|
    (((in_do&_net_2))?sg_in89:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in106:8'b0)|
    (((in_do&_net_2))?data_in105:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in105:8'b0)|
    (((in_do&_net_2))?data_in106:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in107:8'b0)|
    (((in_do&_net_2))?data_in104:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in90:8'b0)|
    (((in_do&_net_2))?data_in89:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b01101010:8'b0)|
    (((in_do&_net_2))?8'b01101001:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_39_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 136 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 89 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_39_add_exe)
  begin
#1 if (_add_map_x_39_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_39_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 136 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 89 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_39_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_39_p_reset = p_reset;
   assign  _add_map_x_39_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in103:128'b0)|
    (((in_do&_net_2))?all_sg_in104:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in105:128'b0)|
    (((in_do&_net_2))?all_sg_in102:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in88:128'b0)|
    (((in_do&_net_2))?all_sg_in87:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)|
    (((in_do&_net_2))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org103:8'b0)|
    (((in_do&_net_2))?data_in_org104:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org105:8'b0)|
    (((in_do&_net_2))?data_in_org102:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org88:8'b0)|
    (((in_do&_net_2))?data_in_org87:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org104:8'b0)|
    (((in_do&_net_2))?data_in_org103:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in103:2'b0)|
    (((in_do&_net_2))?sg_in104:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in105:2'b0)|
    (((in_do&_net_2))?sg_in102:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?2'b00:2'b0)|
    (((in_do&_net_2))?2'b00:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in88:2'b0)|
    (((in_do&_net_2))?sg_in87:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in104:8'b0)|
    (((in_do&_net_2))?data_in103:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in103:8'b0)|
    (((in_do&_net_2))?data_in104:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in105:8'b0)|
    (((in_do&_net_2))?data_in102:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in88:8'b0)|
    (((in_do&_net_2))?data_in87:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b01101000:8'b0)|
    (((in_do&_net_2))?8'b01100111:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_38_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 135 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 88 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_38_add_exe)
  begin
#1 if (_add_map_x_38_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_38_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 135 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 88 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_38_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_38_p_reset = p_reset;
   assign  _add_map_x_38_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in101:128'b0)|
    (((in_do&_net_2))?all_sg_in102:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in103:128'b0)|
    (((in_do&_net_2))?all_sg_in100:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in86:128'b0)|
    (((in_do&_net_2))?all_sg_in85:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)|
    (((in_do&_net_2))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org101:8'b0)|
    (((in_do&_net_2))?data_in_org102:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org103:8'b0)|
    (((in_do&_net_2))?data_in_org100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org86:8'b0)|
    (((in_do&_net_2))?data_in_org85:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org102:8'b0)|
    (((in_do&_net_2))?data_in_org101:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in101:2'b0)|
    (((in_do&_net_2))?sg_in102:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in103:2'b0)|
    (((in_do&_net_2))?sg_in100:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?2'b00:2'b0)|
    (((in_do&_net_2))?2'b00:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in86:2'b0)|
    (((in_do&_net_2))?sg_in85:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in102:8'b0)|
    (((in_do&_net_2))?data_in101:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in101:8'b0)|
    (((in_do&_net_2))?data_in102:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in103:8'b0)|
    (((in_do&_net_2))?data_in100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in86:8'b0)|
    (((in_do&_net_2))?data_in85:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b01100110:8'b0)|
    (((in_do&_net_2))?8'b01100101:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_37_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 134 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 87 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_37_add_exe)
  begin
#1 if (_add_map_x_37_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_37_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 134 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 87 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_37_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_37_p_reset = p_reset;
   assign  _add_map_x_37_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in99:128'b0)|
    (((in_do&_net_2))?all_sg_in100:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in101:128'b0)|
    (((in_do&_net_2))?all_sg_in98:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in84:128'b0)|
    (((in_do&_net_2))?all_sg_in83:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)|
    (((in_do&_net_2))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org99:8'b0)|
    (((in_do&_net_2))?data_in_org100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org101:8'b0)|
    (((in_do&_net_2))?data_in_org98:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org84:8'b0)|
    (((in_do&_net_2))?data_in_org83:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org100:8'b0)|
    (((in_do&_net_2))?data_in_org99:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in99:2'b0)|
    (((in_do&_net_2))?sg_in100:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in101:2'b0)|
    (((in_do&_net_2))?sg_in98:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?2'b00:2'b0)|
    (((in_do&_net_2))?2'b00:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in84:2'b0)|
    (((in_do&_net_2))?sg_in83:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in100:8'b0)|
    (((in_do&_net_2))?data_in99:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in99:8'b0)|
    (((in_do&_net_2))?data_in100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in101:8'b0)|
    (((in_do&_net_2))?data_in98:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in84:8'b0)|
    (((in_do&_net_2))?data_in83:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b01100100:8'b0)|
    (((in_do&_net_2))?8'b01100011:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_36_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 133 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 86 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_36_add_exe)
  begin
#1 if (_add_map_x_36_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_36_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 133 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 86 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_36_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_36_p_reset = p_reset;
   assign  _add_map_x_36_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in97:128'b0)|
    (((in_do&_net_2))?all_sg_in98:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in99:128'b0)|
    (((in_do&_net_2))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in82:128'b0)|
    (((in_do&_net_2))?all_sg_in81:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)|
    (((in_do&_net_2))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org97:8'b0)|
    (((in_do&_net_2))?data_in_org98:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org99:8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org82:8'b0)|
    (((in_do&_net_2))?data_in_org81:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org98:8'b0)|
    (((in_do&_net_2))?data_in_org97:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in97:2'b0)|
    (((in_do&_net_2))?sg_in98:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in99:2'b0)|
    (((in_do&_net_2))?2'b00:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?2'b00:2'b0)|
    (((in_do&_net_2))?2'b00:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in82:2'b0)|
    (((in_do&_net_2))?sg_in81:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in98:8'b0)|
    (((in_do&_net_2))?data_in97:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in97:8'b0)|
    (((in_do&_net_2))?data_in98:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in99:8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in82:8'b0)|
    (((in_do&_net_2))?data_in81:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b01100010:8'b0)|
    (((in_do&_net_2))?8'b01100001:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_35_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 132 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 85 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_35_add_exe)
  begin
#1 if (_add_map_x_35_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_35_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 132 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 85 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_35_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_35_p_reset = p_reset;
   assign  _add_map_x_35_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in109:128'b0)|
    (((in_do&_net_2))?all_sg_in93:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in94:128'b0)|
    (((in_do&_net_2))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in92:128'b0)|
    (((in_do&_net_2))?all_sg_in78:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in77:128'b0)|
    (((in_do&_net_2))?all_sg_in110:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org94:8'b0)|
    (((in_do&_net_2))?data_in_org93:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org92:8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org77:8'b0)|
    (((in_do&_net_2))?data_in_org78:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org109:8'b0)|
    (((in_do&_net_2))?data_in_org110:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org93:8'b0)|
    (((in_do&_net_2))?data_in_org94:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in94:2'b0)|
    (((in_do&_net_2))?sg_in93:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in77:2'b0)|
    (((in_do&_net_2))?2'b00:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in109:2'b0)|
    (((in_do&_net_2))?sg_in110:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in92:2'b0)|
    (((in_do&_net_2))?sg_in78:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in93:8'b0)|
    (((in_do&_net_2))?data_in94:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in94:8'b0)|
    (((in_do&_net_2))?data_in93:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in92:8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in77:8'b0)|
    (((in_do&_net_2))?data_in78:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in109:8'b0)|
    (((in_do&_net_2))?data_in110:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b01011101:8'b0)|
    (((in_do&_net_2))?8'b01011110:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_34_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 131 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 84 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_34_add_exe)
  begin
#1 if (_add_map_x_34_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_34_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 131 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 84 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_34_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_34_p_reset = p_reset;
   assign  _add_map_x_34_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in107:128'b0)|
    (((in_do&_net_2))?all_sg_in91:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in92:128'b0)|
    (((in_do&_net_2))?all_sg_in93:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in90:128'b0)|
    (((in_do&_net_2))?all_sg_in76:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in75:128'b0)|
    (((in_do&_net_2))?all_sg_in108:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org92:8'b0)|
    (((in_do&_net_2))?data_in_org91:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org90:8'b0)|
    (((in_do&_net_2))?data_in_org93:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org75:8'b0)|
    (((in_do&_net_2))?data_in_org76:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org107:8'b0)|
    (((in_do&_net_2))?data_in_org108:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org91:8'b0)|
    (((in_do&_net_2))?data_in_org92:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in92:2'b0)|
    (((in_do&_net_2))?sg_in91:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in75:2'b0)|
    (((in_do&_net_2))?sg_in93:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in107:2'b0)|
    (((in_do&_net_2))?sg_in108:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in90:2'b0)|
    (((in_do&_net_2))?sg_in76:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in91:8'b0)|
    (((in_do&_net_2))?data_in92:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in92:8'b0)|
    (((in_do&_net_2))?data_in91:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in90:8'b0)|
    (((in_do&_net_2))?data_in93:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in75:8'b0)|
    (((in_do&_net_2))?data_in76:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in107:8'b0)|
    (((in_do&_net_2))?data_in108:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b01011011:8'b0)|
    (((in_do&_net_2))?8'b01011100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_33_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 130 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 83 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_33_add_exe)
  begin
#1 if (_add_map_x_33_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_33_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 130 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 83 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_33_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_33_p_reset = p_reset;
   assign  _add_map_x_33_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in105:128'b0)|
    (((in_do&_net_2))?all_sg_in89:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in90:128'b0)|
    (((in_do&_net_2))?all_sg_in91:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in88:128'b0)|
    (((in_do&_net_2))?all_sg_in74:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in73:128'b0)|
    (((in_do&_net_2))?all_sg_in106:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org90:8'b0)|
    (((in_do&_net_2))?data_in_org89:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org88:8'b0)|
    (((in_do&_net_2))?data_in_org91:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org73:8'b0)|
    (((in_do&_net_2))?data_in_org74:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org105:8'b0)|
    (((in_do&_net_2))?data_in_org106:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org89:8'b0)|
    (((in_do&_net_2))?data_in_org90:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in90:2'b0)|
    (((in_do&_net_2))?sg_in89:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in73:2'b0)|
    (((in_do&_net_2))?sg_in91:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in105:2'b0)|
    (((in_do&_net_2))?sg_in106:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in88:2'b0)|
    (((in_do&_net_2))?sg_in74:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in89:8'b0)|
    (((in_do&_net_2))?data_in90:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in90:8'b0)|
    (((in_do&_net_2))?data_in89:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in88:8'b0)|
    (((in_do&_net_2))?data_in91:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in73:8'b0)|
    (((in_do&_net_2))?data_in74:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in105:8'b0)|
    (((in_do&_net_2))?data_in106:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b01011001:8'b0)|
    (((in_do&_net_2))?8'b01011010:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_32_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 129 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 82 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_32_add_exe)
  begin
#1 if (_add_map_x_32_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_32_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 129 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 82 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_32_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_32_p_reset = p_reset;
   assign  _add_map_x_32_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in103:128'b0)|
    (((in_do&_net_2))?all_sg_in87:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in88:128'b0)|
    (((in_do&_net_2))?all_sg_in89:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in86:128'b0)|
    (((in_do&_net_2))?all_sg_in72:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in71:128'b0)|
    (((in_do&_net_2))?all_sg_in104:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org88:8'b0)|
    (((in_do&_net_2))?data_in_org87:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org86:8'b0)|
    (((in_do&_net_2))?data_in_org89:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org71:8'b0)|
    (((in_do&_net_2))?data_in_org72:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org103:8'b0)|
    (((in_do&_net_2))?data_in_org104:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org87:8'b0)|
    (((in_do&_net_2))?data_in_org88:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in88:2'b0)|
    (((in_do&_net_2))?sg_in87:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in71:2'b0)|
    (((in_do&_net_2))?sg_in89:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in103:2'b0)|
    (((in_do&_net_2))?sg_in104:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in86:2'b0)|
    (((in_do&_net_2))?sg_in72:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in87:8'b0)|
    (((in_do&_net_2))?data_in88:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in88:8'b0)|
    (((in_do&_net_2))?data_in87:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in86:8'b0)|
    (((in_do&_net_2))?data_in89:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in71:8'b0)|
    (((in_do&_net_2))?data_in72:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in103:8'b0)|
    (((in_do&_net_2))?data_in104:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b01010111:8'b0)|
    (((in_do&_net_2))?8'b01011000:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_31_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 128 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 81 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_31_add_exe)
  begin
#1 if (_add_map_x_31_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_31_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 128 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 81 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_31_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_31_p_reset = p_reset;
   assign  _add_map_x_31_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in101:128'b0)|
    (((in_do&_net_2))?all_sg_in85:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in86:128'b0)|
    (((in_do&_net_2))?all_sg_in87:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in84:128'b0)|
    (((in_do&_net_2))?all_sg_in70:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in69:128'b0)|
    (((in_do&_net_2))?all_sg_in102:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org86:8'b0)|
    (((in_do&_net_2))?data_in_org85:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org84:8'b0)|
    (((in_do&_net_2))?data_in_org87:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org69:8'b0)|
    (((in_do&_net_2))?data_in_org70:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org101:8'b0)|
    (((in_do&_net_2))?data_in_org102:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org85:8'b0)|
    (((in_do&_net_2))?data_in_org86:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in86:2'b0)|
    (((in_do&_net_2))?sg_in85:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in69:2'b0)|
    (((in_do&_net_2))?sg_in87:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in101:2'b0)|
    (((in_do&_net_2))?sg_in102:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in84:2'b0)|
    (((in_do&_net_2))?sg_in70:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in85:8'b0)|
    (((in_do&_net_2))?data_in86:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in86:8'b0)|
    (((in_do&_net_2))?data_in85:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in84:8'b0)|
    (((in_do&_net_2))?data_in87:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in69:8'b0)|
    (((in_do&_net_2))?data_in70:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in101:8'b0)|
    (((in_do&_net_2))?data_in102:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b01010101:8'b0)|
    (((in_do&_net_2))?8'b01010110:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_30_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 127 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 80 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_30_add_exe)
  begin
#1 if (_add_map_x_30_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_30_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 127 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 80 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_30_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_30_p_reset = p_reset;
   assign  _add_map_x_30_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in99:128'b0)|
    (((in_do&_net_2))?all_sg_in83:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in84:128'b0)|
    (((in_do&_net_2))?all_sg_in85:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in82:128'b0)|
    (((in_do&_net_2))?all_sg_in68:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in67:128'b0)|
    (((in_do&_net_2))?all_sg_in100:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org84:8'b0)|
    (((in_do&_net_2))?data_in_org83:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org82:8'b0)|
    (((in_do&_net_2))?data_in_org85:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org67:8'b0)|
    (((in_do&_net_2))?data_in_org68:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org99:8'b0)|
    (((in_do&_net_2))?data_in_org100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org83:8'b0)|
    (((in_do&_net_2))?data_in_org84:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in84:2'b0)|
    (((in_do&_net_2))?sg_in83:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in67:2'b0)|
    (((in_do&_net_2))?sg_in85:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in99:2'b0)|
    (((in_do&_net_2))?sg_in100:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in82:2'b0)|
    (((in_do&_net_2))?sg_in68:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in83:8'b0)|
    (((in_do&_net_2))?data_in84:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in84:8'b0)|
    (((in_do&_net_2))?data_in83:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in82:8'b0)|
    (((in_do&_net_2))?data_in85:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in67:8'b0)|
    (((in_do&_net_2))?data_in68:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in99:8'b0)|
    (((in_do&_net_2))?data_in100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b01010011:8'b0)|
    (((in_do&_net_2))?8'b01010100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_29_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 126 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 79 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_29_add_exe)
  begin
#1 if (_add_map_x_29_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_29_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 126 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 79 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_29_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_29_p_reset = p_reset;
   assign  _add_map_x_29_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in97:128'b0)|
    (((in_do&_net_2))?all_sg_in81:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in82:128'b0)|
    (((in_do&_net_2))?all_sg_in83:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)|
    (((in_do&_net_2))?all_sg_in66:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in65:128'b0)|
    (((in_do&_net_2))?all_sg_in98:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org82:8'b0)|
    (((in_do&_net_2))?data_in_org81:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?data_in_org83:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org65:8'b0)|
    (((in_do&_net_2))?data_in_org66:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org97:8'b0)|
    (((in_do&_net_2))?data_in_org98:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org81:8'b0)|
    (((in_do&_net_2))?data_in_org82:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in82:2'b0)|
    (((in_do&_net_2))?sg_in81:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in65:2'b0)|
    (((in_do&_net_2))?sg_in83:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in97:2'b0)|
    (((in_do&_net_2))?sg_in98:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?2'b00:2'b0)|
    (((in_do&_net_2))?sg_in66:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in81:8'b0)|
    (((in_do&_net_2))?data_in82:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in82:8'b0)|
    (((in_do&_net_2))?data_in81:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?data_in83:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in65:8'b0)|
    (((in_do&_net_2))?data_in66:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in97:8'b0)|
    (((in_do&_net_2))?data_in98:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b01010001:8'b0)|
    (((in_do&_net_2))?8'b01010010:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_28_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 125 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 78 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_28_add_exe)
  begin
#1 if (_add_map_x_28_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_28_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 125 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 78 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_28_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_28_p_reset = p_reset;
   assign  _add_map_x_28_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in77:128'b0)|
    (((in_do&_net_2))?all_sg_in78:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)|
    (((in_do&_net_2))?all_sg_in76:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in62:128'b0)|
    (((in_do&_net_2))?all_sg_in61:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in94:128'b0)|
    (((in_do&_net_2))?all_sg_in93:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org77:8'b0)|
    (((in_do&_net_2))?data_in_org78:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?data_in_org76:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org62:8'b0)|
    (((in_do&_net_2))?data_in_org61:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org94:8'b0)|
    (((in_do&_net_2))?data_in_org93:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org78:8'b0)|
    (((in_do&_net_2))?data_in_org77:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in77:2'b0)|
    (((in_do&_net_2))?sg_in78:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?2'b00:2'b0)|
    (((in_do&_net_2))?sg_in76:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in94:2'b0)|
    (((in_do&_net_2))?sg_in93:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in62:2'b0)|
    (((in_do&_net_2))?sg_in61:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in78:8'b0)|
    (((in_do&_net_2))?data_in77:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in77:8'b0)|
    (((in_do&_net_2))?data_in78:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?data_in76:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in62:8'b0)|
    (((in_do&_net_2))?data_in61:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in94:8'b0)|
    (((in_do&_net_2))?data_in93:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b01001110:8'b0)|
    (((in_do&_net_2))?8'b01001101:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_27_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 124 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 77 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_27_add_exe)
  begin
#1 if (_add_map_x_27_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_27_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 124 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 77 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_27_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_27_p_reset = p_reset;
   assign  _add_map_x_27_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in75:128'b0)|
    (((in_do&_net_2))?all_sg_in76:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in77:128'b0)|
    (((in_do&_net_2))?all_sg_in74:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in60:128'b0)|
    (((in_do&_net_2))?all_sg_in59:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in92:128'b0)|
    (((in_do&_net_2))?all_sg_in91:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org75:8'b0)|
    (((in_do&_net_2))?data_in_org76:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org77:8'b0)|
    (((in_do&_net_2))?data_in_org74:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org60:8'b0)|
    (((in_do&_net_2))?data_in_org59:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org92:8'b0)|
    (((in_do&_net_2))?data_in_org91:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org76:8'b0)|
    (((in_do&_net_2))?data_in_org75:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in75:2'b0)|
    (((in_do&_net_2))?sg_in76:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in77:2'b0)|
    (((in_do&_net_2))?sg_in74:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in92:2'b0)|
    (((in_do&_net_2))?sg_in91:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in60:2'b0)|
    (((in_do&_net_2))?sg_in59:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in76:8'b0)|
    (((in_do&_net_2))?data_in75:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in75:8'b0)|
    (((in_do&_net_2))?data_in76:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in77:8'b0)|
    (((in_do&_net_2))?data_in74:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in60:8'b0)|
    (((in_do&_net_2))?data_in59:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in92:8'b0)|
    (((in_do&_net_2))?data_in91:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b01001100:8'b0)|
    (((in_do&_net_2))?8'b01001011:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_26_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 123 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 76 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_26_add_exe)
  begin
#1 if (_add_map_x_26_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_26_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 123 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 76 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_26_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_26_p_reset = p_reset;
   assign  _add_map_x_26_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in73:128'b0)|
    (((in_do&_net_2))?all_sg_in74:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in75:128'b0)|
    (((in_do&_net_2))?all_sg_in72:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in58:128'b0)|
    (((in_do&_net_2))?all_sg_in57:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in90:128'b0)|
    (((in_do&_net_2))?all_sg_in89:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org73:8'b0)|
    (((in_do&_net_2))?data_in_org74:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org75:8'b0)|
    (((in_do&_net_2))?data_in_org72:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org58:8'b0)|
    (((in_do&_net_2))?data_in_org57:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org90:8'b0)|
    (((in_do&_net_2))?data_in_org89:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org74:8'b0)|
    (((in_do&_net_2))?data_in_org73:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in73:2'b0)|
    (((in_do&_net_2))?sg_in74:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in75:2'b0)|
    (((in_do&_net_2))?sg_in72:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in90:2'b0)|
    (((in_do&_net_2))?sg_in89:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in58:2'b0)|
    (((in_do&_net_2))?sg_in57:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in74:8'b0)|
    (((in_do&_net_2))?data_in73:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in73:8'b0)|
    (((in_do&_net_2))?data_in74:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in75:8'b0)|
    (((in_do&_net_2))?data_in72:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in58:8'b0)|
    (((in_do&_net_2))?data_in57:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in90:8'b0)|
    (((in_do&_net_2))?data_in89:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b01001010:8'b0)|
    (((in_do&_net_2))?8'b01001001:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_25_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 122 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 75 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_25_add_exe)
  begin
#1 if (_add_map_x_25_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_25_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 122 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 75 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_25_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_25_p_reset = p_reset;
   assign  _add_map_x_25_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in71:128'b0)|
    (((in_do&_net_2))?all_sg_in72:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in73:128'b0)|
    (((in_do&_net_2))?all_sg_in70:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in56:128'b0)|
    (((in_do&_net_2))?all_sg_in55:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in88:128'b0)|
    (((in_do&_net_2))?all_sg_in87:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org71:8'b0)|
    (((in_do&_net_2))?data_in_org72:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org73:8'b0)|
    (((in_do&_net_2))?data_in_org70:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org56:8'b0)|
    (((in_do&_net_2))?data_in_org55:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org88:8'b0)|
    (((in_do&_net_2))?data_in_org87:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org72:8'b0)|
    (((in_do&_net_2))?data_in_org71:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in71:2'b0)|
    (((in_do&_net_2))?sg_in72:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in73:2'b0)|
    (((in_do&_net_2))?sg_in70:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in88:2'b0)|
    (((in_do&_net_2))?sg_in87:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in56:2'b0)|
    (((in_do&_net_2))?sg_in55:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in72:8'b0)|
    (((in_do&_net_2))?data_in71:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in71:8'b0)|
    (((in_do&_net_2))?data_in72:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in73:8'b0)|
    (((in_do&_net_2))?data_in70:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in56:8'b0)|
    (((in_do&_net_2))?data_in55:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in88:8'b0)|
    (((in_do&_net_2))?data_in87:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b01001000:8'b0)|
    (((in_do&_net_2))?8'b01000111:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_24_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 121 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 74 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_24_add_exe)
  begin
#1 if (_add_map_x_24_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_24_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 121 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 74 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_24_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_24_p_reset = p_reset;
   assign  _add_map_x_24_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in69:128'b0)|
    (((in_do&_net_2))?all_sg_in70:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in71:128'b0)|
    (((in_do&_net_2))?all_sg_in68:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in54:128'b0)|
    (((in_do&_net_2))?all_sg_in53:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in86:128'b0)|
    (((in_do&_net_2))?all_sg_in85:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org69:8'b0)|
    (((in_do&_net_2))?data_in_org70:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org71:8'b0)|
    (((in_do&_net_2))?data_in_org68:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org54:8'b0)|
    (((in_do&_net_2))?data_in_org53:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org86:8'b0)|
    (((in_do&_net_2))?data_in_org85:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org70:8'b0)|
    (((in_do&_net_2))?data_in_org69:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in69:2'b0)|
    (((in_do&_net_2))?sg_in70:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in71:2'b0)|
    (((in_do&_net_2))?sg_in68:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in86:2'b0)|
    (((in_do&_net_2))?sg_in85:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in54:2'b0)|
    (((in_do&_net_2))?sg_in53:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in70:8'b0)|
    (((in_do&_net_2))?data_in69:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in69:8'b0)|
    (((in_do&_net_2))?data_in70:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in71:8'b0)|
    (((in_do&_net_2))?data_in68:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in54:8'b0)|
    (((in_do&_net_2))?data_in53:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in86:8'b0)|
    (((in_do&_net_2))?data_in85:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b01000110:8'b0)|
    (((in_do&_net_2))?8'b01000101:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_23_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 120 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 73 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_23_add_exe)
  begin
#1 if (_add_map_x_23_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_23_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 120 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 73 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_23_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_23_p_reset = p_reset;
   assign  _add_map_x_23_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in67:128'b0)|
    (((in_do&_net_2))?all_sg_in68:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in69:128'b0)|
    (((in_do&_net_2))?all_sg_in66:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in52:128'b0)|
    (((in_do&_net_2))?all_sg_in51:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in84:128'b0)|
    (((in_do&_net_2))?all_sg_in83:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org67:8'b0)|
    (((in_do&_net_2))?data_in_org68:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org69:8'b0)|
    (((in_do&_net_2))?data_in_org66:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org52:8'b0)|
    (((in_do&_net_2))?data_in_org51:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org84:8'b0)|
    (((in_do&_net_2))?data_in_org83:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org68:8'b0)|
    (((in_do&_net_2))?data_in_org67:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in67:2'b0)|
    (((in_do&_net_2))?sg_in68:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in69:2'b0)|
    (((in_do&_net_2))?sg_in66:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in84:2'b0)|
    (((in_do&_net_2))?sg_in83:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in52:2'b0)|
    (((in_do&_net_2))?sg_in51:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in68:8'b0)|
    (((in_do&_net_2))?data_in67:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in67:8'b0)|
    (((in_do&_net_2))?data_in68:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in69:8'b0)|
    (((in_do&_net_2))?data_in66:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in52:8'b0)|
    (((in_do&_net_2))?data_in51:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in84:8'b0)|
    (((in_do&_net_2))?data_in83:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b01000100:8'b0)|
    (((in_do&_net_2))?8'b01000011:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_22_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 119 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 72 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_22_add_exe)
  begin
#1 if (_add_map_x_22_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_22_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 119 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 72 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_22_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_22_p_reset = p_reset;
   assign  _add_map_x_22_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in65:128'b0)|
    (((in_do&_net_2))?all_sg_in66:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in67:128'b0)|
    (((in_do&_net_2))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in50:128'b0)|
    (((in_do&_net_2))?all_sg_in49:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in82:128'b0)|
    (((in_do&_net_2))?all_sg_in81:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org65:8'b0)|
    (((in_do&_net_2))?data_in_org66:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org67:8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org50:8'b0)|
    (((in_do&_net_2))?data_in_org49:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org82:8'b0)|
    (((in_do&_net_2))?data_in_org81:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org66:8'b0)|
    (((in_do&_net_2))?data_in_org65:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in65:2'b0)|
    (((in_do&_net_2))?sg_in66:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in67:2'b0)|
    (((in_do&_net_2))?2'b00:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in82:2'b0)|
    (((in_do&_net_2))?sg_in81:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in50:2'b0)|
    (((in_do&_net_2))?sg_in49:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in66:8'b0)|
    (((in_do&_net_2))?data_in65:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in65:8'b0)|
    (((in_do&_net_2))?data_in66:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in67:8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in50:8'b0)|
    (((in_do&_net_2))?data_in49:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in82:8'b0)|
    (((in_do&_net_2))?data_in81:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b01000010:8'b0)|
    (((in_do&_net_2))?8'b01000001:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_21_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 118 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 71 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_21_add_exe)
  begin
#1 if (_add_map_x_21_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_21_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 118 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 71 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_21_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_21_p_reset = p_reset;
   assign  _add_map_x_21_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in77:128'b0)|
    (((in_do&_net_2))?all_sg_in61:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in62:128'b0)|
    (((in_do&_net_2))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in60:128'b0)|
    (((in_do&_net_2))?all_sg_in46:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in45:128'b0)|
    (((in_do&_net_2))?all_sg_in78:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org62:8'b0)|
    (((in_do&_net_2))?data_in_org61:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org60:8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org45:8'b0)|
    (((in_do&_net_2))?data_in_org46:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org77:8'b0)|
    (((in_do&_net_2))?data_in_org78:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org61:8'b0)|
    (((in_do&_net_2))?data_in_org62:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in62:2'b0)|
    (((in_do&_net_2))?sg_in61:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in45:2'b0)|
    (((in_do&_net_2))?2'b00:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in77:2'b0)|
    (((in_do&_net_2))?sg_in78:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in60:2'b0)|
    (((in_do&_net_2))?sg_in46:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in61:8'b0)|
    (((in_do&_net_2))?data_in62:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in62:8'b0)|
    (((in_do&_net_2))?data_in61:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in60:8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in45:8'b0)|
    (((in_do&_net_2))?data_in46:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in77:8'b0)|
    (((in_do&_net_2))?data_in78:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b00111101:8'b0)|
    (((in_do&_net_2))?8'b00111110:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_20_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 117 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 70 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_20_add_exe)
  begin
#1 if (_add_map_x_20_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_20_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 117 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 70 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_20_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_20_p_reset = p_reset;
   assign  _add_map_x_20_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in75:128'b0)|
    (((in_do&_net_2))?all_sg_in59:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in60:128'b0)|
    (((in_do&_net_2))?all_sg_in61:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in58:128'b0)|
    (((in_do&_net_2))?all_sg_in44:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in43:128'b0)|
    (((in_do&_net_2))?all_sg_in76:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org60:8'b0)|
    (((in_do&_net_2))?data_in_org59:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org58:8'b0)|
    (((in_do&_net_2))?data_in_org61:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org43:8'b0)|
    (((in_do&_net_2))?data_in_org44:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org75:8'b0)|
    (((in_do&_net_2))?data_in_org76:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org59:8'b0)|
    (((in_do&_net_2))?data_in_org60:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in60:2'b0)|
    (((in_do&_net_2))?sg_in59:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in43:2'b0)|
    (((in_do&_net_2))?sg_in61:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in75:2'b0)|
    (((in_do&_net_2))?sg_in76:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in58:2'b0)|
    (((in_do&_net_2))?sg_in44:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in59:8'b0)|
    (((in_do&_net_2))?data_in60:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in60:8'b0)|
    (((in_do&_net_2))?data_in59:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in58:8'b0)|
    (((in_do&_net_2))?data_in61:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in43:8'b0)|
    (((in_do&_net_2))?data_in44:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in75:8'b0)|
    (((in_do&_net_2))?data_in76:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b00111011:8'b0)|
    (((in_do&_net_2))?8'b00111100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_19_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 116 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 69 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_19_add_exe)
  begin
#1 if (_add_map_x_19_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_19_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 116 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 69 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_19_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_19_p_reset = p_reset;
   assign  _add_map_x_19_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in73:128'b0)|
    (((in_do&_net_2))?all_sg_in57:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in58:128'b0)|
    (((in_do&_net_2))?all_sg_in59:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in56:128'b0)|
    (((in_do&_net_2))?all_sg_in42:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in41:128'b0)|
    (((in_do&_net_2))?all_sg_in74:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org58:8'b0)|
    (((in_do&_net_2))?data_in_org57:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org56:8'b0)|
    (((in_do&_net_2))?data_in_org59:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org41:8'b0)|
    (((in_do&_net_2))?data_in_org42:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org73:8'b0)|
    (((in_do&_net_2))?data_in_org74:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org57:8'b0)|
    (((in_do&_net_2))?data_in_org58:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in58:2'b0)|
    (((in_do&_net_2))?sg_in57:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in41:2'b0)|
    (((in_do&_net_2))?sg_in59:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in73:2'b0)|
    (((in_do&_net_2))?sg_in74:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in56:2'b0)|
    (((in_do&_net_2))?sg_in42:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in57:8'b0)|
    (((in_do&_net_2))?data_in58:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in58:8'b0)|
    (((in_do&_net_2))?data_in57:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in56:8'b0)|
    (((in_do&_net_2))?data_in59:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in41:8'b0)|
    (((in_do&_net_2))?data_in42:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in73:8'b0)|
    (((in_do&_net_2))?data_in74:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b00111001:8'b0)|
    (((in_do&_net_2))?8'b00111010:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_18_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 115 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 68 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_18_add_exe)
  begin
#1 if (_add_map_x_18_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_18_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 115 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 68 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_18_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_18_p_reset = p_reset;
   assign  _add_map_x_18_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in71:128'b0)|
    (((in_do&_net_2))?all_sg_in55:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in56:128'b0)|
    (((in_do&_net_2))?all_sg_in57:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in54:128'b0)|
    (((in_do&_net_2))?all_sg_in40:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in39:128'b0)|
    (((in_do&_net_2))?all_sg_in72:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org56:8'b0)|
    (((in_do&_net_2))?data_in_org55:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org54:8'b0)|
    (((in_do&_net_2))?data_in_org57:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org39:8'b0)|
    (((in_do&_net_2))?data_in_org40:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org71:8'b0)|
    (((in_do&_net_2))?data_in_org72:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org55:8'b0)|
    (((in_do&_net_2))?data_in_org56:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in56:2'b0)|
    (((in_do&_net_2))?sg_in55:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in39:2'b0)|
    (((in_do&_net_2))?sg_in57:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in71:2'b0)|
    (((in_do&_net_2))?sg_in72:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in54:2'b0)|
    (((in_do&_net_2))?sg_in40:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in55:8'b0)|
    (((in_do&_net_2))?data_in56:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in56:8'b0)|
    (((in_do&_net_2))?data_in55:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in54:8'b0)|
    (((in_do&_net_2))?data_in57:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in39:8'b0)|
    (((in_do&_net_2))?data_in40:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in71:8'b0)|
    (((in_do&_net_2))?data_in72:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b00110111:8'b0)|
    (((in_do&_net_2))?8'b00111000:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_17_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 114 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 67 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_17_add_exe)
  begin
#1 if (_add_map_x_17_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_17_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 114 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 67 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_17_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_17_p_reset = p_reset;
   assign  _add_map_x_17_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in69:128'b0)|
    (((in_do&_net_2))?all_sg_in53:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in54:128'b0)|
    (((in_do&_net_2))?all_sg_in55:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in52:128'b0)|
    (((in_do&_net_2))?all_sg_in38:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in37:128'b0)|
    (((in_do&_net_2))?all_sg_in70:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org54:8'b0)|
    (((in_do&_net_2))?data_in_org53:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org52:8'b0)|
    (((in_do&_net_2))?data_in_org55:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org37:8'b0)|
    (((in_do&_net_2))?data_in_org38:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org69:8'b0)|
    (((in_do&_net_2))?data_in_org70:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org53:8'b0)|
    (((in_do&_net_2))?data_in_org54:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in54:2'b0)|
    (((in_do&_net_2))?sg_in53:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in37:2'b0)|
    (((in_do&_net_2))?sg_in55:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in69:2'b0)|
    (((in_do&_net_2))?sg_in70:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in52:2'b0)|
    (((in_do&_net_2))?sg_in38:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in53:8'b0)|
    (((in_do&_net_2))?data_in54:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in54:8'b0)|
    (((in_do&_net_2))?data_in53:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in52:8'b0)|
    (((in_do&_net_2))?data_in55:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in37:8'b0)|
    (((in_do&_net_2))?data_in38:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in69:8'b0)|
    (((in_do&_net_2))?data_in70:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b00110101:8'b0)|
    (((in_do&_net_2))?8'b00110110:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_16_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 113 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 66 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_16_add_exe)
  begin
#1 if (_add_map_x_16_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_16_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 113 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 66 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_16_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_16_p_reset = p_reset;
   assign  _add_map_x_16_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in67:128'b0)|
    (((in_do&_net_2))?all_sg_in51:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in52:128'b0)|
    (((in_do&_net_2))?all_sg_in53:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in50:128'b0)|
    (((in_do&_net_2))?all_sg_in36:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in35:128'b0)|
    (((in_do&_net_2))?all_sg_in68:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org52:8'b0)|
    (((in_do&_net_2))?data_in_org51:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org50:8'b0)|
    (((in_do&_net_2))?data_in_org53:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org35:8'b0)|
    (((in_do&_net_2))?data_in_org36:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org67:8'b0)|
    (((in_do&_net_2))?data_in_org68:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org51:8'b0)|
    (((in_do&_net_2))?data_in_org52:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in52:2'b0)|
    (((in_do&_net_2))?sg_in51:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in35:2'b0)|
    (((in_do&_net_2))?sg_in53:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in67:2'b0)|
    (((in_do&_net_2))?sg_in68:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in50:2'b0)|
    (((in_do&_net_2))?sg_in36:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in51:8'b0)|
    (((in_do&_net_2))?data_in52:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in52:8'b0)|
    (((in_do&_net_2))?data_in51:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in50:8'b0)|
    (((in_do&_net_2))?data_in53:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in35:8'b0)|
    (((in_do&_net_2))?data_in36:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in67:8'b0)|
    (((in_do&_net_2))?data_in68:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b00110011:8'b0)|
    (((in_do&_net_2))?8'b00110100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_15_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 112 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 65 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_15_add_exe)
  begin
#1 if (_add_map_x_15_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_15_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 112 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 65 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_15_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_15_p_reset = p_reset;
   assign  _add_map_x_15_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in65:128'b0)|
    (((in_do&_net_2))?all_sg_in49:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in50:128'b0)|
    (((in_do&_net_2))?all_sg_in51:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)|
    (((in_do&_net_2))?all_sg_in34:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in33:128'b0)|
    (((in_do&_net_2))?all_sg_in66:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org50:8'b0)|
    (((in_do&_net_2))?data_in_org49:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?data_in_org51:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org33:8'b0)|
    (((in_do&_net_2))?data_in_org34:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org65:8'b0)|
    (((in_do&_net_2))?data_in_org66:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org49:8'b0)|
    (((in_do&_net_2))?data_in_org50:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in50:2'b0)|
    (((in_do&_net_2))?sg_in49:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in33:2'b0)|
    (((in_do&_net_2))?sg_in51:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in65:2'b0)|
    (((in_do&_net_2))?sg_in66:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?2'b00:2'b0)|
    (((in_do&_net_2))?sg_in34:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in49:8'b0)|
    (((in_do&_net_2))?data_in50:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in50:8'b0)|
    (((in_do&_net_2))?data_in49:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?data_in51:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in33:8'b0)|
    (((in_do&_net_2))?data_in34:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in65:8'b0)|
    (((in_do&_net_2))?data_in66:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b00110001:8'b0)|
    (((in_do&_net_2))?8'b00110010:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_14_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 111 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 64 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_14_add_exe)
  begin
#1 if (_add_map_x_14_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_14_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 111 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 64 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_14_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_14_p_reset = p_reset;
   assign  _add_map_x_14_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in45:128'b0)|
    (((in_do&_net_2))?all_sg_in46:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)|
    (((in_do&_net_2))?all_sg_in44:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in30:128'b0)|
    (((in_do&_net_2))?all_sg_in29:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in62:128'b0)|
    (((in_do&_net_2))?all_sg_in61:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org45:8'b0)|
    (((in_do&_net_2))?data_in_org46:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?data_in_org44:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org30:8'b0)|
    (((in_do&_net_2))?data_in_org29:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org62:8'b0)|
    (((in_do&_net_2))?data_in_org61:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org46:8'b0)|
    (((in_do&_net_2))?data_in_org45:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in45:2'b0)|
    (((in_do&_net_2))?sg_in46:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?2'b00:2'b0)|
    (((in_do&_net_2))?sg_in44:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in62:2'b0)|
    (((in_do&_net_2))?sg_in61:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in30:2'b0)|
    (((in_do&_net_2))?sg_in29:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in46:8'b0)|
    (((in_do&_net_2))?data_in45:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in45:8'b0)|
    (((in_do&_net_2))?data_in46:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?data_in44:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in30:8'b0)|
    (((in_do&_net_2))?data_in29:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in62:8'b0)|
    (((in_do&_net_2))?data_in61:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b00101110:8'b0)|
    (((in_do&_net_2))?8'b00101101:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_13_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 110 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 63 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_13_add_exe)
  begin
#1 if (_add_map_x_13_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_13_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 110 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 63 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_13_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_13_p_reset = p_reset;
   assign  _add_map_x_13_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in43:128'b0)|
    (((in_do&_net_2))?all_sg_in44:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in45:128'b0)|
    (((in_do&_net_2))?all_sg_in42:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in28:128'b0)|
    (((in_do&_net_2))?all_sg_in27:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in60:128'b0)|
    (((in_do&_net_2))?all_sg_in59:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org43:8'b0)|
    (((in_do&_net_2))?data_in_org44:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org45:8'b0)|
    (((in_do&_net_2))?data_in_org42:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org28:8'b0)|
    (((in_do&_net_2))?data_in_org27:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org60:8'b0)|
    (((in_do&_net_2))?data_in_org59:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org44:8'b0)|
    (((in_do&_net_2))?data_in_org43:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in43:2'b0)|
    (((in_do&_net_2))?sg_in44:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in45:2'b0)|
    (((in_do&_net_2))?sg_in42:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in60:2'b0)|
    (((in_do&_net_2))?sg_in59:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in28:2'b0)|
    (((in_do&_net_2))?sg_in27:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in44:8'b0)|
    (((in_do&_net_2))?data_in43:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in43:8'b0)|
    (((in_do&_net_2))?data_in44:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in45:8'b0)|
    (((in_do&_net_2))?data_in42:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in28:8'b0)|
    (((in_do&_net_2))?data_in27:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in60:8'b0)|
    (((in_do&_net_2))?data_in59:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b00101100:8'b0)|
    (((in_do&_net_2))?8'b00101011:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_12_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 109 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 62 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_12_add_exe)
  begin
#1 if (_add_map_x_12_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_12_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 109 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 62 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_12_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_12_p_reset = p_reset;
   assign  _add_map_x_12_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in41:128'b0)|
    (((in_do&_net_2))?all_sg_in42:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in43:128'b0)|
    (((in_do&_net_2))?all_sg_in40:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in26:128'b0)|
    (((in_do&_net_2))?all_sg_in25:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in58:128'b0)|
    (((in_do&_net_2))?all_sg_in57:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org41:8'b0)|
    (((in_do&_net_2))?data_in_org42:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org43:8'b0)|
    (((in_do&_net_2))?data_in_org40:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org26:8'b0)|
    (((in_do&_net_2))?data_in_org25:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org58:8'b0)|
    (((in_do&_net_2))?data_in_org57:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org42:8'b0)|
    (((in_do&_net_2))?data_in_org41:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in41:2'b0)|
    (((in_do&_net_2))?sg_in42:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in43:2'b0)|
    (((in_do&_net_2))?sg_in40:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in58:2'b0)|
    (((in_do&_net_2))?sg_in57:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in26:2'b0)|
    (((in_do&_net_2))?sg_in25:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in42:8'b0)|
    (((in_do&_net_2))?data_in41:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in41:8'b0)|
    (((in_do&_net_2))?data_in42:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in43:8'b0)|
    (((in_do&_net_2))?data_in40:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in26:8'b0)|
    (((in_do&_net_2))?data_in25:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in58:8'b0)|
    (((in_do&_net_2))?data_in57:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b00101010:8'b0)|
    (((in_do&_net_2))?8'b00101001:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_11_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 108 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 61 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_11_add_exe)
  begin
#1 if (_add_map_x_11_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_11_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 108 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 61 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_11_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_11_p_reset = p_reset;
   assign  _add_map_x_11_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in39:128'b0)|
    (((in_do&_net_2))?all_sg_in40:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in41:128'b0)|
    (((in_do&_net_2))?all_sg_in38:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in24:128'b0)|
    (((in_do&_net_2))?all_sg_in23:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in56:128'b0)|
    (((in_do&_net_2))?all_sg_in55:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org39:8'b0)|
    (((in_do&_net_2))?data_in_org40:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org41:8'b0)|
    (((in_do&_net_2))?data_in_org38:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org24:8'b0)|
    (((in_do&_net_2))?data_in_org23:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org56:8'b0)|
    (((in_do&_net_2))?data_in_org55:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org40:8'b0)|
    (((in_do&_net_2))?data_in_org39:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in39:2'b0)|
    (((in_do&_net_2))?sg_in40:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in41:2'b0)|
    (((in_do&_net_2))?sg_in38:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in56:2'b0)|
    (((in_do&_net_2))?sg_in55:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in24:2'b0)|
    (((in_do&_net_2))?sg_in23:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in40:8'b0)|
    (((in_do&_net_2))?data_in39:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in39:8'b0)|
    (((in_do&_net_2))?data_in40:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in41:8'b0)|
    (((in_do&_net_2))?data_in38:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in24:8'b0)|
    (((in_do&_net_2))?data_in23:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in56:8'b0)|
    (((in_do&_net_2))?data_in55:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b00101000:8'b0)|
    (((in_do&_net_2))?8'b00100111:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_10_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 107 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 60 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_10_add_exe)
  begin
#1 if (_add_map_x_10_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_10_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 107 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 60 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_10_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_10_p_reset = p_reset;
   assign  _add_map_x_10_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in37:128'b0)|
    (((in_do&_net_2))?all_sg_in38:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in39:128'b0)|
    (((in_do&_net_2))?all_sg_in36:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in22:128'b0)|
    (((in_do&_net_2))?all_sg_in21:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in54:128'b0)|
    (((in_do&_net_2))?all_sg_in53:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org37:8'b0)|
    (((in_do&_net_2))?data_in_org38:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org39:8'b0)|
    (((in_do&_net_2))?data_in_org36:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org22:8'b0)|
    (((in_do&_net_2))?data_in_org21:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org54:8'b0)|
    (((in_do&_net_2))?data_in_org53:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org38:8'b0)|
    (((in_do&_net_2))?data_in_org37:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in37:2'b0)|
    (((in_do&_net_2))?sg_in38:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in39:2'b0)|
    (((in_do&_net_2))?sg_in36:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in54:2'b0)|
    (((in_do&_net_2))?sg_in53:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in22:2'b0)|
    (((in_do&_net_2))?sg_in21:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in38:8'b0)|
    (((in_do&_net_2))?data_in37:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in37:8'b0)|
    (((in_do&_net_2))?data_in38:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in39:8'b0)|
    (((in_do&_net_2))?data_in36:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in22:8'b0)|
    (((in_do&_net_2))?data_in21:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in54:8'b0)|
    (((in_do&_net_2))?data_in53:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b00100110:8'b0)|
    (((in_do&_net_2))?8'b00100101:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_9_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 106 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 59 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_9_add_exe)
  begin
#1 if (_add_map_x_9_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_9_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 106 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 59 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_9_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_9_p_reset = p_reset;
   assign  _add_map_x_9_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in35:128'b0)|
    (((in_do&_net_2))?all_sg_in36:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in37:128'b0)|
    (((in_do&_net_2))?all_sg_in34:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in20:128'b0)|
    (((in_do&_net_2))?all_sg_in19:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in52:128'b0)|
    (((in_do&_net_2))?all_sg_in51:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org35:8'b0)|
    (((in_do&_net_2))?data_in_org36:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org37:8'b0)|
    (((in_do&_net_2))?data_in_org34:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org20:8'b0)|
    (((in_do&_net_2))?data_in_org19:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org52:8'b0)|
    (((in_do&_net_2))?data_in_org51:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org36:8'b0)|
    (((in_do&_net_2))?data_in_org35:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in35:2'b0)|
    (((in_do&_net_2))?sg_in36:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in37:2'b0)|
    (((in_do&_net_2))?sg_in34:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in52:2'b0)|
    (((in_do&_net_2))?sg_in51:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in20:2'b0)|
    (((in_do&_net_2))?sg_in19:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in36:8'b0)|
    (((in_do&_net_2))?data_in35:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in35:8'b0)|
    (((in_do&_net_2))?data_in36:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in37:8'b0)|
    (((in_do&_net_2))?data_in34:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in20:8'b0)|
    (((in_do&_net_2))?data_in19:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in52:8'b0)|
    (((in_do&_net_2))?data_in51:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b00100100:8'b0)|
    (((in_do&_net_2))?8'b00100011:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_8_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 105 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 58 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_8_add_exe)
  begin
#1 if (_add_map_x_8_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_8_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 105 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 58 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_8_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_8_p_reset = p_reset;
   assign  _add_map_x_8_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in33:128'b0)|
    (((in_do&_net_2))?all_sg_in34:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in35:128'b0)|
    (((in_do&_net_2))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in18:128'b0)|
    (((in_do&_net_2))?all_sg_in17:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in50:128'b0)|
    (((in_do&_net_2))?all_sg_in49:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org33:8'b0)|
    (((in_do&_net_2))?data_in_org34:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org35:8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org18:8'b0)|
    (((in_do&_net_2))?data_in_org17:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org50:8'b0)|
    (((in_do&_net_2))?data_in_org49:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org34:8'b0)|
    (((in_do&_net_2))?data_in_org33:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in33:2'b0)|
    (((in_do&_net_2))?sg_in34:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in35:2'b0)|
    (((in_do&_net_2))?2'b00:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in50:2'b0)|
    (((in_do&_net_2))?sg_in49:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in18:2'b0)|
    (((in_do&_net_2))?sg_in17:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in34:8'b0)|
    (((in_do&_net_2))?data_in33:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in33:8'b0)|
    (((in_do&_net_2))?data_in34:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in35:8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in18:8'b0)|
    (((in_do&_net_2))?data_in17:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in50:8'b0)|
    (((in_do&_net_2))?data_in49:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b00100010:8'b0)|
    (((in_do&_net_2))?8'b00100001:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_7_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 104 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 57 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_7_add_exe)
  begin
#1 if (_add_map_x_7_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_7_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 104 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 57 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_7_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_7_p_reset = p_reset;
   assign  _add_map_x_7_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in45:128'b0)|
    (((in_do&_net_2))?all_sg_in29:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in30:128'b0)|
    (((in_do&_net_2))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in28:128'b0)|
    (((in_do&_net_2))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)|
    (((in_do&_net_2))?all_sg_in46:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org30:8'b0)|
    (((in_do&_net_2))?data_in_org29:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org28:8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org45:8'b0)|
    (((in_do&_net_2))?data_in_org46:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org29:8'b0)|
    (((in_do&_net_2))?data_in_org30:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in30:2'b0)|
    (((in_do&_net_2))?sg_in29:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?2'b00:2'b0)|
    (((in_do&_net_2))?2'b00:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in45:2'b0)|
    (((in_do&_net_2))?sg_in46:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in28:2'b0)|
    (((in_do&_net_2))?2'b00:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in29:8'b0)|
    (((in_do&_net_2))?data_in30:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in30:8'b0)|
    (((in_do&_net_2))?data_in29:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in28:8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in45:8'b0)|
    (((in_do&_net_2))?data_in46:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b00011101:8'b0)|
    (((in_do&_net_2))?8'b00011110:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_6_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 103 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 56 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_6_add_exe)
  begin
#1 if (_add_map_x_6_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_6_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 103 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 56 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_6_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_6_p_reset = p_reset;
   assign  _add_map_x_6_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in43:128'b0)|
    (((in_do&_net_2))?all_sg_in27:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in28:128'b0)|
    (((in_do&_net_2))?all_sg_in29:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in26:128'b0)|
    (((in_do&_net_2))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)|
    (((in_do&_net_2))?all_sg_in44:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org28:8'b0)|
    (((in_do&_net_2))?data_in_org27:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org26:8'b0)|
    (((in_do&_net_2))?data_in_org29:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org43:8'b0)|
    (((in_do&_net_2))?data_in_org44:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org27:8'b0)|
    (((in_do&_net_2))?data_in_org28:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in28:2'b0)|
    (((in_do&_net_2))?sg_in27:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?2'b00:2'b0)|
    (((in_do&_net_2))?sg_in29:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in43:2'b0)|
    (((in_do&_net_2))?sg_in44:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in26:2'b0)|
    (((in_do&_net_2))?2'b00:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in27:8'b0)|
    (((in_do&_net_2))?data_in28:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in28:8'b0)|
    (((in_do&_net_2))?data_in27:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in26:8'b0)|
    (((in_do&_net_2))?data_in29:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in43:8'b0)|
    (((in_do&_net_2))?data_in44:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b00011011:8'b0)|
    (((in_do&_net_2))?8'b00011100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_5_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 102 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 55 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_5_add_exe)
  begin
#1 if (_add_map_x_5_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_5_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 102 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 55 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_5_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_5_p_reset = p_reset;
   assign  _add_map_x_5_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in41:128'b0)|
    (((in_do&_net_2))?all_sg_in25:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in26:128'b0)|
    (((in_do&_net_2))?all_sg_in27:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in24:128'b0)|
    (((in_do&_net_2))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)|
    (((in_do&_net_2))?all_sg_in42:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org26:8'b0)|
    (((in_do&_net_2))?data_in_org25:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org24:8'b0)|
    (((in_do&_net_2))?data_in_org27:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org41:8'b0)|
    (((in_do&_net_2))?data_in_org42:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org25:8'b0)|
    (((in_do&_net_2))?data_in_org26:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in26:2'b0)|
    (((in_do&_net_2))?sg_in25:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?2'b00:2'b0)|
    (((in_do&_net_2))?sg_in27:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in41:2'b0)|
    (((in_do&_net_2))?sg_in42:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in24:2'b0)|
    (((in_do&_net_2))?2'b00:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in25:8'b0)|
    (((in_do&_net_2))?data_in26:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in26:8'b0)|
    (((in_do&_net_2))?data_in25:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in24:8'b0)|
    (((in_do&_net_2))?data_in27:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in41:8'b0)|
    (((in_do&_net_2))?data_in42:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b00011001:8'b0)|
    (((in_do&_net_2))?8'b00011010:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_4_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 101 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 54 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_4_add_exe)
  begin
#1 if (_add_map_x_4_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_4_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 101 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 54 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_4_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_4_p_reset = p_reset;
   assign  _add_map_x_4_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in39:128'b0)|
    (((in_do&_net_2))?all_sg_in23:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in24:128'b0)|
    (((in_do&_net_2))?all_sg_in25:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in22:128'b0)|
    (((in_do&_net_2))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)|
    (((in_do&_net_2))?all_sg_in40:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org24:8'b0)|
    (((in_do&_net_2))?data_in_org23:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org22:8'b0)|
    (((in_do&_net_2))?data_in_org25:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org39:8'b0)|
    (((in_do&_net_2))?data_in_org40:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org23:8'b0)|
    (((in_do&_net_2))?data_in_org24:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in24:2'b0)|
    (((in_do&_net_2))?sg_in23:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?2'b00:2'b0)|
    (((in_do&_net_2))?sg_in25:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in39:2'b0)|
    (((in_do&_net_2))?sg_in40:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in22:2'b0)|
    (((in_do&_net_2))?2'b00:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in23:8'b0)|
    (((in_do&_net_2))?data_in24:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in24:8'b0)|
    (((in_do&_net_2))?data_in23:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in22:8'b0)|
    (((in_do&_net_2))?data_in25:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in39:8'b0)|
    (((in_do&_net_2))?data_in40:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b00010111:8'b0)|
    (((in_do&_net_2))?8'b00011000:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_3_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 100 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 53 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_3_add_exe)
  begin
#1 if (_add_map_x_3_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_3_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 100 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 53 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_3_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_3_p_reset = p_reset;
   assign  _add_map_x_3_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in37:128'b0)|
    (((in_do&_net_2))?all_sg_in21:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in22:128'b0)|
    (((in_do&_net_2))?all_sg_in23:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in20:128'b0)|
    (((in_do&_net_2))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)|
    (((in_do&_net_2))?all_sg_in38:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org22:8'b0)|
    (((in_do&_net_2))?data_in_org21:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org20:8'b0)|
    (((in_do&_net_2))?data_in_org23:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org37:8'b0)|
    (((in_do&_net_2))?data_in_org38:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org21:8'b0)|
    (((in_do&_net_2))?data_in_org22:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in22:2'b0)|
    (((in_do&_net_2))?sg_in21:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?2'b00:2'b0)|
    (((in_do&_net_2))?sg_in23:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in37:2'b0)|
    (((in_do&_net_2))?sg_in38:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in20:2'b0)|
    (((in_do&_net_2))?2'b00:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in21:8'b0)|
    (((in_do&_net_2))?data_in22:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in22:8'b0)|
    (((in_do&_net_2))?data_in21:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in20:8'b0)|
    (((in_do&_net_2))?data_in23:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in37:8'b0)|
    (((in_do&_net_2))?data_in38:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b00010101:8'b0)|
    (((in_do&_net_2))?8'b00010110:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_2_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 99 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 52 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_2_add_exe)
  begin
#1 if (_add_map_x_2_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_2_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 99 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 52 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_2_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_2_p_reset = p_reset;
   assign  _add_map_x_2_m_clock = m_clock;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_wall_end_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_wall_end_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?wall_end_in:128'b0)|
    (((in_do&_net_2))?wall_end_in:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_all_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_all_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in35:128'b0)|
    (((in_do&_net_2))?all_sg_in19:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_all_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_all_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in20:128'b0)|
    (((in_do&_net_2))?all_sg_in21:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_all_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_all_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?all_sg_in18:128'b0)|
    (((in_do&_net_2))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_all_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_all_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 128'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000:128'b0)|
    (((in_do&_net_2))?all_sg_in36:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_moto_org_near) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_moto_org_near = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org20:8'b0)|
    (((in_do&_net_2))?data_in_org19:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_moto_org_near1) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_moto_org_near1 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org18:8'b0)|
    (((in_do&_net_2))?data_in_org21:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_moto_org_near2) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_moto_org_near2 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_moto_org_near3) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_moto_org_near3 = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org35:8'b0)|
    (((in_do&_net_2))?data_in_org36:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_moto_org) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_moto_org = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in_org19:8'b0)|
    (((in_do&_net_2))?data_in_org20:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_sg_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_sg_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in20:2'b0)|
    (((in_do&_net_2))?sg_in19:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_sg_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_sg_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?2'b00:2'b0)|
    (((in_do&_net_2))?sg_in21:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_sg_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_sg_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in35:2'b0)|
    (((in_do&_net_2))?sg_in36:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_sg_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_sg_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 2'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?sg_in18:2'b0)|
    (((in_do&_net_2))?2'b00:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_wall_t_in) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_wall_t_in = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 1'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?dig_w:1'b0)|
    (((in_do&_net_2))?dig_w:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_moto) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_moto = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in19:8'b0)|
    (((in_do&_net_2))?data_in20:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_up) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_up = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in20:8'b0)|
    (((in_do&_net_2))?data_in19:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_right) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_right = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in18:8'b0)|
    (((in_do&_net_2))?data_in21:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_down) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_down = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)|
    (((in_do&_net_2))?({({1'b1,1'b1,1'b1,1'b1,1'b1,1'b1,1'b1}),1'b1}):8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_left) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_left = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?data_in35:8'b0)|
    (((in_do&_net_2))?data_in36:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_start) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_start = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?start:8'b0)|
    (((in_do&_net_2))?start:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_goal) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_goal = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?goal:8'b0)|
    (((in_do&_net_2))?goal:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_now) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_now = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?8'b00010011:8'b0)|
    (((in_do&_net_2))?8'b00010100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if (((in_do&_net_3)&(in_do&_net_2)))
 begin $display("Warning: assign collision(add_all:_add_map_x_1_distance) at %d",$time);
if ((in_do&_net_3)) $display("assert ((in_do&_net_3)) line 98 at %d\n",$time);
if ((in_do&_net_2)) $display("assert ((in_do&_net_2)) line 51 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_distance = 
// synthesis translate_off
// synopsys translate_off
(((in_do&_net_3)&(in_do&_net_2)))? 8'bx :(((in_do&_net_3)|(in_do&_net_2)))? 
// synthesis translate_on
// synopsys translate_on
(((in_do&_net_3))?distance_count_all:8'b0)|
    (((in_do&_net_2))?distance_count_all:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _add_map_x_1_add_exe)
  begin
#1 if (_add_map_x_1_add_exe===1'bx)
 begin
$display("Warning: control hazard(add_all:_add_map_x_1_add_exe) at %d",$time);
 end
#1 if ((((in_do&_net_3))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_3) || 1'b1) line 98 at %d\n",$time);
#1 if ((((in_do&_net_2))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do&_net_2) || 1'b1) line 51 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _add_map_x_1_add_exe = (in_do&_net_3)|
    (in_do&_net_2);
   assign  _add_map_x_1_p_reset = p_reset;
   assign  _add_map_x_1_m_clock = m_clock;
   assign  _net_0 = (sig_reg==1'b1);
   assign  _net_1 = (sig_reg==1'b0);
   assign  _net_2 = 
// synthesis translate_off
// synopsys translate_off
(in_do)? 
// synthesis translate_on
// synopsys translate_on
((in_do)?(sig==1'b1):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _net_3 = 
// synthesis translate_off
// synopsys translate_off
(in_do)? 
// synthesis translate_on
// synopsys translate_on
((in_do)?(sig==1'b0):1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t0) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t0 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t1) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t1 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_1_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_1_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t2) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t2 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_2_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_2_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t3) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t3 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_3_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_3_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t4) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t4 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_4_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_4_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t5) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t5 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_5_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_5_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t6) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t6 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_6_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_6_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t7) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t7 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_7_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_7_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t8) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t8 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_8_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_8_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t9) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t9 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_9_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_9_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t10) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t10 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_10_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_10_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t11) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t11 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_11_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_11_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t12) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t12 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_12_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_12_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t13) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t13 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_13_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_13_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t14) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t14 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_14_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_14_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t15) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t15 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_15_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_15_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t16) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t16 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_16_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_16_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t17) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t17 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_17_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_17_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t18) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t18 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_18_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_18_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t19) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t19 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_19_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_19_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t20) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t20 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_20_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_20_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t21) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t21 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_21_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_21_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t22) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t22 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_22_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_22_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t23) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t23 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_23_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_23_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t24) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t24 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_24_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_24_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t25) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t25 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_25_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_25_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t26) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t26 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_26_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_26_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t27) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t27 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_27_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_27_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t28) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t28 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_28_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_28_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t29) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t29 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_29_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_29_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t30) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t30 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_30_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_30_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t31) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t31 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_31_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_31_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t32) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t32 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_32_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_32_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t33) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t33 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_33_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_33_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t34) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t34 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_34_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_34_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t35) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t35 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_35_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_35_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t36) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t36 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_36_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_36_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t37) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t37 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_37_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_37_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t38) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t38 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_38_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_38_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t39) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t39 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_39_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_39_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t40) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t40 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_40_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_40_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:dig_t41) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  dig_t41 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 1'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_41_wall_t_out:1'b0)|
    ((_net_0)?_add_map_x_41_wall_t_out:1'b0)
// synthesis translate_off
// synopsys translate_off
:1'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:wall_end) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  wall_end = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?(((((((((((((((((((((((((((((((((((((((((_add_map_x_end_wall|_add_map_x_1_end_wall)|_add_map_x_2_end_wall)|_add_map_x_3_end_wall)|_add_map_x_4_end_wall)|_add_map_x_5_end_wall)|_add_map_x_6_end_wall)|_add_map_x_7_end_wall)|_add_map_x_8_end_wall)|_add_map_x_9_end_wall)|_add_map_x_10_end_wall)|_add_map_x_11_end_wall)|_add_map_x_12_end_wall)|_add_map_x_13_end_wall)|_add_map_x_14_end_wall)|_add_map_x_15_end_wall)|_add_map_x_16_end_wall)|_add_map_x_17_end_wall)|_add_map_x_18_end_wall)|_add_map_x_19_end_wall)|_add_map_x_20_end_wall)|_add_map_x_21_end_wall)|_add_map_x_22_end_wall)|_add_map_x_23_end_wall)|_add_map_x_24_end_wall)|_add_map_x_25_end_wall)|_add_map_x_26_end_wall)|_add_map_x_27_end_wall)|_add_map_x_28_end_wall)|_add_map_x_29_end_wall)|_add_map_x_30_end_wall)|_add_map_x_31_end_wall)|_add_map_x_32_end_wall)|_add_map_x_33_end_wall)|_add_map_x_34_end_wall)|_add_map_x_35_end_wall)|_add_map_x_36_end_wall)|_add_map_x_37_end_wall)|_add_map_x_38_end_wall)|_add_map_x_39_end_wall)|_add_map_x_40_end_wall)|_add_map_x_41_end_wall):128'b0)|
    ((_net_0)?(((((((((((((((((((((((((((((((((((((((((_add_map_x_end_wall|_add_map_x_1_end_wall)|_add_map_x_2_end_wall)|_add_map_x_3_end_wall)|_add_map_x_4_end_wall)|_add_map_x_5_end_wall)|_add_map_x_6_end_wall)|_add_map_x_7_end_wall)|_add_map_x_8_end_wall)|_add_map_x_9_end_wall)|_add_map_x_10_end_wall)|_add_map_x_11_end_wall)|_add_map_x_12_end_wall)|_add_map_x_13_end_wall)|_add_map_x_14_end_wall)|_add_map_x_15_end_wall)|_add_map_x_16_end_wall)|_add_map_x_17_end_wall)|_add_map_x_18_end_wall)|_add_map_x_19_end_wall)|_add_map_x_20_end_wall)|_add_map_x_21_end_wall)|_add_map_x_22_end_wall)|_add_map_x_23_end_wall)|_add_map_x_24_end_wall)|_add_map_x_25_end_wall)|_add_map_x_26_end_wall)|_add_map_x_27_end_wall)|_add_map_x_28_end_wall)|_add_map_x_29_end_wall)|_add_map_x_30_end_wall)|_add_map_x_31_end_wall)|_add_map_x_32_end_wall)|_add_map_x_33_end_wall)|_add_map_x_34_end_wall)|_add_map_x_35_end_wall)|_add_map_x_36_end_wall)|_add_map_x_37_end_wall)|_add_map_x_38_end_wall)|_add_map_x_39_end_wall)|_add_map_x_40_end_wall)|_add_map_x_41_end_wall):128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org17) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org17 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_data_org:8'b0)|
    ((_net_0)?_add_map_x_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org18) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org18 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org19) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org19 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_1_data_org:8'b0)|
    ((_net_0)?_add_map_x_1_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org20) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org20 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_1_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_1_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org21) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org21 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_2_data_org:8'b0)|
    ((_net_0)?_add_map_x_2_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org22) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org22 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_2_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_2_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org23) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org23 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_3_data_org:8'b0)|
    ((_net_0)?_add_map_x_3_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org24) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org24 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_3_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_3_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org25) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org25 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_4_data_org:8'b0)|
    ((_net_0)?_add_map_x_4_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org26) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org26 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_4_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_4_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org27) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org27 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_5_data_org:8'b0)|
    ((_net_0)?_add_map_x_5_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org28) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org28 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_5_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_5_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org29) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org29 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_6_data_org:8'b0)|
    ((_net_0)?_add_map_x_6_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org30) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org30 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_6_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_6_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org33) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org33 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_7_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_7_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org34) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org34 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_7_data_org:8'b0)|
    ((_net_0)?_add_map_x_7_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org35) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org35 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_8_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_8_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org36) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org36 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_8_data_org:8'b0)|
    ((_net_0)?_add_map_x_8_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org37) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org37 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_9_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_9_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org38) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org38 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_9_data_org:8'b0)|
    ((_net_0)?_add_map_x_9_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org39) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org39 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_10_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_10_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org40) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org40 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_10_data_org:8'b0)|
    ((_net_0)?_add_map_x_10_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org41) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org41 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_11_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_11_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org42) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org42 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_11_data_org:8'b0)|
    ((_net_0)?_add_map_x_11_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org43) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org43 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_12_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_12_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org44) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org44 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_12_data_org:8'b0)|
    ((_net_0)?_add_map_x_12_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org45) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org45 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_13_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_13_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org46) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org46 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_13_data_org:8'b0)|
    ((_net_0)?_add_map_x_13_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org49) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org49 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_14_data_org:8'b0)|
    ((_net_0)?_add_map_x_14_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org50) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org50 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_14_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_14_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org51) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org51 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_15_data_org:8'b0)|
    ((_net_0)?_add_map_x_15_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org52) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org52 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_15_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_15_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org53) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org53 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_16_data_org:8'b0)|
    ((_net_0)?_add_map_x_16_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org54) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org54 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_16_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_16_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org55) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org55 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_17_data_org:8'b0)|
    ((_net_0)?_add_map_x_17_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org56) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org56 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_17_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_17_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org57) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org57 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_18_data_org:8'b0)|
    ((_net_0)?_add_map_x_18_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org58) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org58 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_18_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_18_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org59) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org59 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_19_data_org:8'b0)|
    ((_net_0)?_add_map_x_19_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org60) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org60 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_19_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_19_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org61) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org61 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_20_data_org:8'b0)|
    ((_net_0)?_add_map_x_20_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org62) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org62 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_20_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_20_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org65) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org65 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_21_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_21_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org66) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org66 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_21_data_org:8'b0)|
    ((_net_0)?_add_map_x_21_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org67) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org67 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_22_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_22_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org68) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org68 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_22_data_org:8'b0)|
    ((_net_0)?_add_map_x_22_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org69) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org69 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_23_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_23_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org70) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org70 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_23_data_org:8'b0)|
    ((_net_0)?_add_map_x_23_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org71) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org71 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_24_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_24_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org72) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org72 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_24_data_org:8'b0)|
    ((_net_0)?_add_map_x_24_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org73) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org73 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_25_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_25_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org74) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org74 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_25_data_org:8'b0)|
    ((_net_0)?_add_map_x_25_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org75) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org75 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_26_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_26_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org76) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org76 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_26_data_org:8'b0)|
    ((_net_0)?_add_map_x_26_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org77) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org77 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_27_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_27_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org78) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org78 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_27_data_org:8'b0)|
    ((_net_0)?_add_map_x_27_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org81) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org81 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_28_data_org:8'b0)|
    ((_net_0)?_add_map_x_28_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org82) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org82 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_28_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_28_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org83) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org83 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_29_data_org:8'b0)|
    ((_net_0)?_add_map_x_29_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org84) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org84 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_29_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_29_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org85) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org85 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_30_data_org:8'b0)|
    ((_net_0)?_add_map_x_30_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org86) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org86 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_30_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_30_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org87) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org87 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_31_data_org:8'b0)|
    ((_net_0)?_add_map_x_31_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org88) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org88 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_31_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_31_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org89) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org89 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_32_data_org:8'b0)|
    ((_net_0)?_add_map_x_32_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org90) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org90 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_32_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_32_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org91) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org91 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_33_data_org:8'b0)|
    ((_net_0)?_add_map_x_33_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org92) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org92 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_33_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_33_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org93) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org93 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_34_data_org:8'b0)|
    ((_net_0)?_add_map_x_34_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org94) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org94 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_34_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_34_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org97) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org97 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_35_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_35_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org98) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org98 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_35_data_org:8'b0)|
    ((_net_0)?_add_map_x_35_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org99) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org99 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_36_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_36_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org100) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org100 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_36_data_org:8'b0)|
    ((_net_0)?_add_map_x_36_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org101) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org101 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_37_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_37_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org102) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org102 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_37_data_org:8'b0)|
    ((_net_0)?_add_map_x_37_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org103) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org103 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_38_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_38_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org104) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org104 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_38_data_org:8'b0)|
    ((_net_0)?_add_map_x_38_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org105) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org105 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_39_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_39_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org106) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org106 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_39_data_org:8'b0)|
    ((_net_0)?_add_map_x_39_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org107) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org107 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_40_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_40_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org108) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org108 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_40_data_org:8'b0)|
    ((_net_0)?_add_map_x_40_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org109) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org109 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_41_data_org_near:8'b0)|
    ((_net_0)?_add_map_x_41_data_org:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_org110) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_org110 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_41_data_org:8'b0)|
    ((_net_0)?_add_map_x_41_data_org_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out17) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out17 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_s_g:2'b0)|
    ((_net_0)?_add_map_x_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out18) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out18 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out19) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out19 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_1_s_g:2'b0)|
    ((_net_0)?_add_map_x_1_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out20) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out20 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_1_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_1_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out21) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out21 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_2_s_g:2'b0)|
    ((_net_0)?_add_map_x_2_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out22) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out22 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_2_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_2_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out23) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out23 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_3_s_g:2'b0)|
    ((_net_0)?_add_map_x_3_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out24) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out24 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_3_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_3_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out25) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out25 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_4_s_g:2'b0)|
    ((_net_0)?_add_map_x_4_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out26) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out26 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_4_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_4_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out27) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out27 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_5_s_g:2'b0)|
    ((_net_0)?_add_map_x_5_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out28) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out28 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_5_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_5_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out29) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out29 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_6_s_g:2'b0)|
    ((_net_0)?_add_map_x_6_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out30) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out30 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_6_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_6_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out33) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out33 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_7_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_7_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out34) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out34 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_7_s_g:2'b0)|
    ((_net_0)?_add_map_x_7_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out35) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out35 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_8_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_8_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out36) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out36 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_8_s_g:2'b0)|
    ((_net_0)?_add_map_x_8_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out37) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out37 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_9_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_9_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out38) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out38 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_9_s_g:2'b0)|
    ((_net_0)?_add_map_x_9_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out39) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out39 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_10_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_10_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out40) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out40 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_10_s_g:2'b0)|
    ((_net_0)?_add_map_x_10_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out41) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out41 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_11_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_11_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out42) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out42 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_11_s_g:2'b0)|
    ((_net_0)?_add_map_x_11_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out43) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out43 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_12_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_12_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out44) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out44 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_12_s_g:2'b0)|
    ((_net_0)?_add_map_x_12_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out45) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out45 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_13_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_13_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out46) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out46 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_13_s_g:2'b0)|
    ((_net_0)?_add_map_x_13_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out49) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out49 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_14_s_g:2'b0)|
    ((_net_0)?_add_map_x_14_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out50) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out50 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_14_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_14_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out51) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out51 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_15_s_g:2'b0)|
    ((_net_0)?_add_map_x_15_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out52) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out52 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_15_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_15_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out53) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out53 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_16_s_g:2'b0)|
    ((_net_0)?_add_map_x_16_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out54) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out54 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_16_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_16_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out55) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out55 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_17_s_g:2'b0)|
    ((_net_0)?_add_map_x_17_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out56) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out56 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_17_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_17_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out57) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out57 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_18_s_g:2'b0)|
    ((_net_0)?_add_map_x_18_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out58) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out58 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_18_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_18_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out59) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out59 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_19_s_g:2'b0)|
    ((_net_0)?_add_map_x_19_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out60) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out60 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_19_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_19_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out61) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out61 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_20_s_g:2'b0)|
    ((_net_0)?_add_map_x_20_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out62) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out62 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_20_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_20_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out65) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out65 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_21_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_21_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out66) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out66 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_21_s_g:2'b0)|
    ((_net_0)?_add_map_x_21_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out67) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out67 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_22_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_22_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out68) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out68 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_22_s_g:2'b0)|
    ((_net_0)?_add_map_x_22_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out69) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out69 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_23_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_23_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out70) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out70 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_23_s_g:2'b0)|
    ((_net_0)?_add_map_x_23_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out71) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out71 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_24_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_24_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out72) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out72 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_24_s_g:2'b0)|
    ((_net_0)?_add_map_x_24_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out73) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out73 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_25_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_25_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out74) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out74 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_25_s_g:2'b0)|
    ((_net_0)?_add_map_x_25_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out75) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out75 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_26_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_26_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out76) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out76 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_26_s_g:2'b0)|
    ((_net_0)?_add_map_x_26_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out77) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out77 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_27_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_27_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out78) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out78 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_27_s_g:2'b0)|
    ((_net_0)?_add_map_x_27_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out81) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out81 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_28_s_g:2'b0)|
    ((_net_0)?_add_map_x_28_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out82) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out82 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_28_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_28_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out83) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out83 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_29_s_g:2'b0)|
    ((_net_0)?_add_map_x_29_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out84) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out84 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_29_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_29_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out85) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out85 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_30_s_g:2'b0)|
    ((_net_0)?_add_map_x_30_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out86) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out86 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_30_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_30_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out87) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out87 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_31_s_g:2'b0)|
    ((_net_0)?_add_map_x_31_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out88) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out88 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_31_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_31_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out89) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out89 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_32_s_g:2'b0)|
    ((_net_0)?_add_map_x_32_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out90) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out90 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_32_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_32_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out91) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out91 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_33_s_g:2'b0)|
    ((_net_0)?_add_map_x_33_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out92) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out92 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_33_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_33_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out93) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out93 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_34_s_g:2'b0)|
    ((_net_0)?_add_map_x_34_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out94) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out94 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_34_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_34_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out97) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out97 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_35_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_35_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out98) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out98 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_35_s_g:2'b0)|
    ((_net_0)?_add_map_x_35_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out99) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out99 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_36_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_36_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out100) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out100 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_36_s_g:2'b0)|
    ((_net_0)?_add_map_x_36_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out101) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out101 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_37_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_37_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out102) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out102 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_37_s_g:2'b0)|
    ((_net_0)?_add_map_x_37_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out103) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out103 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_38_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_38_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out104) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out104 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_38_s_g:2'b0)|
    ((_net_0)?_add_map_x_38_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out105) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out105 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_39_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_39_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out106) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out106 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_39_s_g:2'b0)|
    ((_net_0)?_add_map_x_39_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out107) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out107 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_40_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_40_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out108) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out108 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_40_s_g:2'b0)|
    ((_net_0)?_add_map_x_40_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out109) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out109 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_41_s_g_near:2'b0)|
    ((_net_0)?_add_map_x_41_s_g:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:sg_out110) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  sg_out110 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 2'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_41_s_g:2'b0)|
    ((_net_0)?_add_map_x_41_s_g_near:2'b0)
// synthesis translate_off
// synopsys translate_off
:2'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out17) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out17 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_data_out:8'b0)|
    ((_net_0)?_add_map_x_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out18) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out18 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_data_near:8'b0)|
    ((_net_0)?_add_map_x_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out19) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out19 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_1_data_out:8'b0)|
    ((_net_0)?_add_map_x_1_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out20) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out20 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_1_data_near:8'b0)|
    ((_net_0)?_add_map_x_1_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out21) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out21 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_2_data_out:8'b0)|
    ((_net_0)?_add_map_x_2_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out22) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out22 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_2_data_near:8'b0)|
    ((_net_0)?_add_map_x_2_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out23) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out23 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_3_data_out:8'b0)|
    ((_net_0)?_add_map_x_3_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out24) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out24 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_3_data_near:8'b0)|
    ((_net_0)?_add_map_x_3_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out25) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out25 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_4_data_out:8'b0)|
    ((_net_0)?_add_map_x_4_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out26) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out26 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_4_data_near:8'b0)|
    ((_net_0)?_add_map_x_4_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out27) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out27 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_5_data_out:8'b0)|
    ((_net_0)?_add_map_x_5_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out28) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out28 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_5_data_near:8'b0)|
    ((_net_0)?_add_map_x_5_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out29) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out29 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_6_data_out:8'b0)|
    ((_net_0)?_add_map_x_6_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out30) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out30 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_6_data_near:8'b0)|
    ((_net_0)?_add_map_x_6_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out33) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out33 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_7_data_near:8'b0)|
    ((_net_0)?_add_map_x_7_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out34) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out34 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_7_data_out:8'b0)|
    ((_net_0)?_add_map_x_7_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out35) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out35 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_8_data_near:8'b0)|
    ((_net_0)?_add_map_x_8_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out36) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out36 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_8_data_out:8'b0)|
    ((_net_0)?_add_map_x_8_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out37) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out37 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_9_data_near:8'b0)|
    ((_net_0)?_add_map_x_9_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out38) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out38 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_9_data_out:8'b0)|
    ((_net_0)?_add_map_x_9_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out39) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out39 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_10_data_near:8'b0)|
    ((_net_0)?_add_map_x_10_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out40) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out40 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_10_data_out:8'b0)|
    ((_net_0)?_add_map_x_10_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out41) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out41 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_11_data_near:8'b0)|
    ((_net_0)?_add_map_x_11_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out42) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out42 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_11_data_out:8'b0)|
    ((_net_0)?_add_map_x_11_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out43) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out43 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_12_data_near:8'b0)|
    ((_net_0)?_add_map_x_12_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out44) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out44 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_12_data_out:8'b0)|
    ((_net_0)?_add_map_x_12_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out45) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out45 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_13_data_near:8'b0)|
    ((_net_0)?_add_map_x_13_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out46) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out46 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_13_data_out:8'b0)|
    ((_net_0)?_add_map_x_13_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out49) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out49 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_14_data_out:8'b0)|
    ((_net_0)?_add_map_x_14_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out50) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out50 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_14_data_near:8'b0)|
    ((_net_0)?_add_map_x_14_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out51) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out51 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_15_data_out:8'b0)|
    ((_net_0)?_add_map_x_15_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out52) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out52 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_15_data_near:8'b0)|
    ((_net_0)?_add_map_x_15_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out53) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out53 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_16_data_out:8'b0)|
    ((_net_0)?_add_map_x_16_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out54) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out54 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_16_data_near:8'b0)|
    ((_net_0)?_add_map_x_16_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out55) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out55 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_17_data_out:8'b0)|
    ((_net_0)?_add_map_x_17_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out56) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out56 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_17_data_near:8'b0)|
    ((_net_0)?_add_map_x_17_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out57) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out57 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_18_data_out:8'b0)|
    ((_net_0)?_add_map_x_18_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out58) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out58 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_18_data_near:8'b0)|
    ((_net_0)?_add_map_x_18_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out59) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out59 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_19_data_out:8'b0)|
    ((_net_0)?_add_map_x_19_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out60) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out60 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_19_data_near:8'b0)|
    ((_net_0)?_add_map_x_19_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out61) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out61 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_20_data_out:8'b0)|
    ((_net_0)?_add_map_x_20_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out62) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out62 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_20_data_near:8'b0)|
    ((_net_0)?_add_map_x_20_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out65) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out65 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_21_data_near:8'b0)|
    ((_net_0)?_add_map_x_21_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out66) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out66 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_21_data_out:8'b0)|
    ((_net_0)?_add_map_x_21_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out67) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out67 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_22_data_near:8'b0)|
    ((_net_0)?_add_map_x_22_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out68) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out68 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_22_data_out:8'b0)|
    ((_net_0)?_add_map_x_22_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out69) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out69 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_23_data_near:8'b0)|
    ((_net_0)?_add_map_x_23_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out70) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out70 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_23_data_out:8'b0)|
    ((_net_0)?_add_map_x_23_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out71) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out71 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_24_data_near:8'b0)|
    ((_net_0)?_add_map_x_24_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out72) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out72 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_24_data_out:8'b0)|
    ((_net_0)?_add_map_x_24_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out73) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out73 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_25_data_near:8'b0)|
    ((_net_0)?_add_map_x_25_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out74) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out74 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_25_data_out:8'b0)|
    ((_net_0)?_add_map_x_25_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out75) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out75 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_26_data_near:8'b0)|
    ((_net_0)?_add_map_x_26_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out76) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out76 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_26_data_out:8'b0)|
    ((_net_0)?_add_map_x_26_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out77) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out77 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_27_data_near:8'b0)|
    ((_net_0)?_add_map_x_27_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out78) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out78 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_27_data_out:8'b0)|
    ((_net_0)?_add_map_x_27_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out81) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out81 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_28_data_out:8'b0)|
    ((_net_0)?_add_map_x_28_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out82) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out82 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_28_data_near:8'b0)|
    ((_net_0)?_add_map_x_28_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out83) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out83 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_29_data_out:8'b0)|
    ((_net_0)?_add_map_x_29_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out84) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out84 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_29_data_near:8'b0)|
    ((_net_0)?_add_map_x_29_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out85) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out85 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_30_data_out:8'b0)|
    ((_net_0)?_add_map_x_30_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out86) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out86 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_30_data_near:8'b0)|
    ((_net_0)?_add_map_x_30_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out87) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out87 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_31_data_out:8'b0)|
    ((_net_0)?_add_map_x_31_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out88) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out88 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_31_data_near:8'b0)|
    ((_net_0)?_add_map_x_31_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out89) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out89 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_32_data_out:8'b0)|
    ((_net_0)?_add_map_x_32_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out90) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out90 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_32_data_near:8'b0)|
    ((_net_0)?_add_map_x_32_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out91) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out91 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_33_data_out:8'b0)|
    ((_net_0)?_add_map_x_33_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out92) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out92 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_33_data_near:8'b0)|
    ((_net_0)?_add_map_x_33_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out93) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out93 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_34_data_out:8'b0)|
    ((_net_0)?_add_map_x_34_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out94) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out94 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_34_data_near:8'b0)|
    ((_net_0)?_add_map_x_34_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out97) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out97 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_35_data_near:8'b0)|
    ((_net_0)?_add_map_x_35_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out98) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out98 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_35_data_out:8'b0)|
    ((_net_0)?_add_map_x_35_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out99) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out99 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_36_data_near:8'b0)|
    ((_net_0)?_add_map_x_36_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out100) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out100 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_36_data_out:8'b0)|
    ((_net_0)?_add_map_x_36_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out101) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out101 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_37_data_near:8'b0)|
    ((_net_0)?_add_map_x_37_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out102) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out102 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_37_data_out:8'b0)|
    ((_net_0)?_add_map_x_37_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out103) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out103 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_38_data_near:8'b0)|
    ((_net_0)?_add_map_x_38_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out104) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out104 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_38_data_out:8'b0)|
    ((_net_0)?_add_map_x_38_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out105) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out105 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_39_data_near:8'b0)|
    ((_net_0)?_add_map_x_39_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out106) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out106 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_39_data_out:8'b0)|
    ((_net_0)?_add_map_x_39_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out107) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out107 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_40_data_near:8'b0)|
    ((_net_0)?_add_map_x_40_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out108) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out108 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_40_data_out:8'b0)|
    ((_net_0)?_add_map_x_40_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out109) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out109 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_41_data_near:8'b0)|
    ((_net_0)?_add_map_x_41_data_out:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out110) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out110 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_41_data_out:8'b0)|
    ((_net_0)?_add_map_x_41_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index17) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index17 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index18) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index18 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_data_near:8'b0)|
    ((_net_0)?_add_map_x_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index19) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index19 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_1_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_1_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index20) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index20 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_1_data_near:8'b0)|
    ((_net_0)?_add_map_x_1_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index21) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index21 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_2_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_2_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index22) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index22 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_2_data_near:8'b0)|
    ((_net_0)?_add_map_x_2_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index23) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index23 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_3_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_3_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index24) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index24 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_3_data_near:8'b0)|
    ((_net_0)?_add_map_x_3_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index25) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index25 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_4_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_4_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index26) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index26 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_4_data_near:8'b0)|
    ((_net_0)?_add_map_x_4_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index27) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index27 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_5_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_5_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index28) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index28 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_5_data_near:8'b0)|
    ((_net_0)?_add_map_x_5_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index29) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index29 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_6_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_6_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index30) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index30 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_6_data_near:8'b0)|
    ((_net_0)?_add_map_x_6_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index33) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index33 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_7_data_near:8'b0)|
    ((_net_0)?_add_map_x_7_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index34) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index34 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_7_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_7_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index35) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index35 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_8_data_near:8'b0)|
    ((_net_0)?_add_map_x_8_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index36) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index36 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_8_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_8_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index37) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index37 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_9_data_near:8'b0)|
    ((_net_0)?_add_map_x_9_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index38) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index38 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_9_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_9_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index39) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index39 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_10_data_near:8'b0)|
    ((_net_0)?_add_map_x_10_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index40) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index40 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_10_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_10_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index41) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index41 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_11_data_near:8'b0)|
    ((_net_0)?_add_map_x_11_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index42) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index42 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_11_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_11_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index43) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index43 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_12_data_near:8'b0)|
    ((_net_0)?_add_map_x_12_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index44) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index44 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_12_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_12_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index45) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index45 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_13_data_near:8'b0)|
    ((_net_0)?_add_map_x_13_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index46) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index46 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_13_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_13_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index49) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index49 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_14_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_14_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index50) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index50 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_14_data_near:8'b0)|
    ((_net_0)?_add_map_x_14_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index51) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index51 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_15_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_15_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index52) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index52 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_15_data_near:8'b0)|
    ((_net_0)?_add_map_x_15_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index53) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index53 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_16_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_16_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index54) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index54 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_16_data_near:8'b0)|
    ((_net_0)?_add_map_x_16_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index55) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index55 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_17_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_17_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index56) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index56 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_17_data_near:8'b0)|
    ((_net_0)?_add_map_x_17_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index57) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index57 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_18_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_18_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index58) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index58 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_18_data_near:8'b0)|
    ((_net_0)?_add_map_x_18_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index59) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index59 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_19_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_19_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index60) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index60 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_19_data_near:8'b0)|
    ((_net_0)?_add_map_x_19_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index61) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index61 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_20_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_20_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index62) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index62 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_20_data_near:8'b0)|
    ((_net_0)?_add_map_x_20_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index65) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index65 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_21_data_near:8'b0)|
    ((_net_0)?_add_map_x_21_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index66) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index66 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_21_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_21_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index67) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index67 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_22_data_near:8'b0)|
    ((_net_0)?_add_map_x_22_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index68) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index68 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_22_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_22_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index69) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index69 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_23_data_near:8'b0)|
    ((_net_0)?_add_map_x_23_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index70) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index70 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_23_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_23_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index71) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index71 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_24_data_near:8'b0)|
    ((_net_0)?_add_map_x_24_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index72) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index72 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_24_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_24_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index73) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index73 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_25_data_near:8'b0)|
    ((_net_0)?_add_map_x_25_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index74) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index74 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_25_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_25_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index75) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index75 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_26_data_near:8'b0)|
    ((_net_0)?_add_map_x_26_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index76) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index76 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_26_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_26_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index77) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index77 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_27_data_near:8'b0)|
    ((_net_0)?_add_map_x_27_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index78) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index78 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_27_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_27_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index81) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index81 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_28_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_28_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index82) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index82 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_28_data_near:8'b0)|
    ((_net_0)?_add_map_x_28_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index83) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index83 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_29_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_29_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index84) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index84 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_29_data_near:8'b0)|
    ((_net_0)?_add_map_x_29_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index85) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index85 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_30_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_30_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index86) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index86 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_30_data_near:8'b0)|
    ((_net_0)?_add_map_x_30_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index87) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index87 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_31_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_31_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index88) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index88 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_31_data_near:8'b0)|
    ((_net_0)?_add_map_x_31_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index89) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index89 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_32_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_32_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index90) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index90 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_32_data_near:8'b0)|
    ((_net_0)?_add_map_x_32_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index91) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index91 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_33_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_33_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index92) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index92 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_33_data_near:8'b0)|
    ((_net_0)?_add_map_x_33_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index93) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index93 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_34_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_34_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index94) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index94 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_34_data_near:8'b0)|
    ((_net_0)?_add_map_x_34_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index97) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index97 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_35_data_near:8'b0)|
    ((_net_0)?_add_map_x_35_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index98) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index98 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_35_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_35_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index99) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index99 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_36_data_near:8'b0)|
    ((_net_0)?_add_map_x_36_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index100) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index100 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_36_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_36_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index101) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index101 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_37_data_near:8'b0)|
    ((_net_0)?_add_map_x_37_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index102) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index102 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_37_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_37_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index103) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index103 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_38_data_near:8'b0)|
    ((_net_0)?_add_map_x_38_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index104) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index104 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_38_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_38_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index105) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index105 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_39_data_near:8'b0)|
    ((_net_0)?_add_map_x_39_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index106) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index106 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_39_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_39_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index107) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index107 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_40_data_near:8'b0)|
    ((_net_0)?_add_map_x_40_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index108) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index108 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_40_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_40_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index109) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index109 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_41_data_near:8'b0)|
    ((_net_0)?_add_map_x_41_data_out_index:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:data_out_index110) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  data_out_index110 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 8'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_41_data_out_index:8'b0)|
    ((_net_0)?_add_map_x_41_data_near:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out17) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out17 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out18) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out18 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out19) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out19 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_1_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_1_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out20) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out20 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_1_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_1_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out21) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out21 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_2_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_2_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out22) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out22 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_2_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_2_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out23) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out23 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_3_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_3_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out24) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out24 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_3_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_3_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out25) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out25 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_4_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_4_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out26) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out26 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_4_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_4_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out27) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out27 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_5_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_5_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out28) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out28 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_5_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_5_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out29) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out29 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_6_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_6_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out30) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out30 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_6_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_6_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out33) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out33 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_7_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_7_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out34) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out34 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_7_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_7_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out35) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out35 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_8_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_8_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out36) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out36 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_8_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_8_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out37) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out37 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_9_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_9_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out38) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out38 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_9_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_9_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out39) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out39 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_10_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_10_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out40) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out40 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_10_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_10_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out41) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out41 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_11_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_11_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out42) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out42 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_11_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_11_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out43) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out43 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_12_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_12_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out44) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out44 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_12_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_12_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out45) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out45 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_13_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_13_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out46) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out46 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_13_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_13_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out49) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out49 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_14_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_14_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out50) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out50 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_14_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_14_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out51) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out51 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_15_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_15_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out52) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out52 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_15_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_15_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out53) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out53 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_16_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_16_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out54) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out54 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_16_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_16_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out55) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out55 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_17_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_17_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out56) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out56 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_17_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_17_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out57) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out57 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_18_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_18_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out58) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out58 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_18_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_18_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out59) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out59 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_19_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_19_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out60) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out60 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_19_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_19_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out61) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out61 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_20_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_20_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out62) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out62 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_20_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_20_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out65) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out65 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_21_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_21_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out66) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out66 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_21_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_21_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out67) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out67 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_22_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_22_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out68) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out68 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_22_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_22_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out69) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out69 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_23_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_23_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out70) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out70 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_23_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_23_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out71) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out71 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_24_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_24_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out72) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out72 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_24_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_24_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out73) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out73 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_25_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_25_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out74) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out74 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_25_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_25_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out75) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out75 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_26_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_26_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out76) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out76 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_26_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_26_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out77) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out77 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_27_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_27_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out78) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out78 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_27_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_27_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out81) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out81 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_28_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_28_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out82) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out82 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_28_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_28_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out83) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out83 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_29_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_29_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out84) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out84 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_29_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_29_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out85) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out85 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_30_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_30_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out86) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out86 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_30_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_30_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out87) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out87 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_31_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_31_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out88) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out88 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_31_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_31_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out89) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out89 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_32_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_32_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out90) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out90 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_32_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_32_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out91) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out91 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_33_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_33_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out92) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out92 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_33_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_33_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out93) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out93 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_34_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_34_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out94) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out94 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_34_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_34_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out97) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out97 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_35_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_35_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out98) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out98 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_35_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_35_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out99) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out99 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_36_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_36_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out100) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out100 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_36_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_36_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out101) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out101 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_37_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_37_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out102) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out102 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_37_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_37_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out103) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out103 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_38_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_38_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out104) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out104 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_38_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_38_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out105) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out105 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_39_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_39_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out106) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out106 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_39_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_39_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out107) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out107 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_40_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_40_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out108) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out108 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_40_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_40_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out109) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out109 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_41_all_s_g_near:128'b0)|
    ((_net_0)?_add_map_x_41_all_s_g:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge m_clock or posedge p_reset)
  begin
if ((_net_1&_net_0))
 begin $display("Warning: assign collision(add_all:all_sg_out110) at %d",$time);
if (_net_1) $display("assert (_net_1) line 38 at %d\n",$time);
if (_net_0) $display("assert (_net_0) line 21 at %d\n",$time);
 end
 end

// synthesis translate_on
// synopsys translate_on
   assign  all_sg_out110 = 
// synthesis translate_off
// synopsys translate_off
((_net_1&_net_0))? 128'bx :((_net_1|_net_0))? 
// synthesis translate_on
// synopsys translate_on
((_net_1)?_add_map_x_41_all_s_g:128'b0)|
    ((_net_0)?_add_map_x_41_all_s_g_near:128'b0)
// synthesis translate_off
// synopsys translate_off
:128'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge out_do)
  begin
#1 if (out_do===1'bx)
 begin
$display("Warning: control hazard(add_all:out_do) at %d",$time);
 end
#1 if (((in_do)===1'bx) || (1'b1)===1'bx) $display("hazard (in_do || 1'b1) line 142 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  out_do = in_do;

// synthesis translate_off
// synopsys translate_off
always @(posedge out_data)
  begin
#1 if (out_data===1'bx)
 begin
$display("Warning: control hazard(add_all:out_data) at %d",$time);
 end
#1 if (((_net_1)===1'bx) || (1'b1)===1'bx) $display("hazard (_net_1 || 1'b1) line 38 at %d\n",$time);
#1 if (((_net_0)===1'bx) || (1'b1)===1'bx) $display("hazard (_net_0 || 1'b1) line 21 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  out_data = _net_1|
    _net_0;
always @(posedge m_clock or posedge p_reset)
  begin
if (p_reset)
     sig_reg <= 1'b0;
else if (in_do)
      sig_reg <= sig;
end
endmodule

/*Produced by NSL Core(version=20240424), IP ARCH, Inc. Tue May 21 04:56:15 2024
 Licensed to :EVALUATION USER*/
