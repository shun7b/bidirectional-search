
/*Produced by NSL Core(version=20240424), IP ARCH, Inc. Tue May 21 04:56:16 2024
 Licensed to :EVALUATION USER*/
/*
 DO NOT USE ANY PART OF THIS FILE FOR COMMERCIAL PRODUCTS. 
*/

module seach ( p_reset , m_clock , data_in17 , data_in18 , data_in19 , data_in20 , data_in21 , data_in22 , data_in23 , data_in24 , data_in25 , data_in26 , data_in27 , data_in28 , data_in29 , data_in30 , data_in33 , data_in34 , data_in35 , data_in36 , data_in37 , data_in38 , data_in39 , data_in40 , data_in41 , data_in42 , data_in43 , data_in44 , data_in45 , data_in46 , data_in49 , data_in50 , data_in51 , data_in52 , data_in53 , data_in54 , data_in55 , data_in56 , data_in57 , data_in58 , data_in59 , data_in60 , data_in61 , data_in62 , data_in65 , data_in66 , data_in67 , data_in68 , data_in69 , data_in70 , data_in71 , data_in72 , data_in73 , data_in74 , data_in75 , data_in76 , data_in77 , data_in78 , data_in81 , data_in82 , data_in83 , data_in84 , data_in85 , data_in86 , data_in87 , data_in88 , data_in89 , data_in90 , data_in91 , data_in92 , data_in93 , data_in94 , data_in97 , data_in98 , data_in99 , data_in100 , data_in101 , data_in102 , data_in103 , data_in104 , data_in105 , data_in106 , data_in107 , data_in108 , data_in109 , data_in110 , data_out17 , data_out18 , data_out19 , data_out20 , data_out21 , data_out22 , data_out23 , data_out24 , data_out25 , data_out26 , data_out27 , data_out28 , data_out29 , data_out30 , data_out33 , data_out34 , data_out35 , data_out36 , data_out37 , data_out38 , data_out39 , data_out40 , data_out41 , data_out42 , data_out43 , data_out44 , data_out45 , data_out46 , data_out49 , data_out50 , data_out51 , data_out52 , data_out53 , data_out54 , data_out55 , data_out56 , data_out57 , data_out58 , data_out59 , data_out60 , data_out61 , data_out62 , data_out65 , data_out66 , data_out67 , data_out68 , data_out69 , data_out70 , data_out71 , data_out72 , data_out73 , data_out74 , data_out75 , data_out76 , data_out77 , data_out78 , data_out81 , data_out82 , data_out83 , data_out84 , data_out85 , data_out86 , data_out87 , data_out88 , data_out89 , data_out90 , data_out91 , data_out92 , data_out93 , data_out94 , data_out97 , data_out98 , data_out99 , data_out100 , data_out101 , data_out102 , data_out103 , data_out104 , data_out105 , data_out106 , data_out107 , data_out108 , data_out109 , data_out110 , startplot , goalplot , in_do , out_do , out_data );
  input p_reset, m_clock;
  wire p_reset, m_clock;
  input [7:0] data_in17;
  wire [7:0] data_in17;
  input [7:0] data_in18;
  wire [7:0] data_in18;
  input [7:0] data_in19;
  wire [7:0] data_in19;
  input [7:0] data_in20;
  wire [7:0] data_in20;
  input [7:0] data_in21;
  wire [7:0] data_in21;
  input [7:0] data_in22;
  wire [7:0] data_in22;
  input [7:0] data_in23;
  wire [7:0] data_in23;
  input [7:0] data_in24;
  wire [7:0] data_in24;
  input [7:0] data_in25;
  wire [7:0] data_in25;
  input [7:0] data_in26;
  wire [7:0] data_in26;
  input [7:0] data_in27;
  wire [7:0] data_in27;
  input [7:0] data_in28;
  wire [7:0] data_in28;
  input [7:0] data_in29;
  wire [7:0] data_in29;
  input [7:0] data_in30;
  wire [7:0] data_in30;
  input [7:0] data_in33;
  wire [7:0] data_in33;
  input [7:0] data_in34;
  wire [7:0] data_in34;
  input [7:0] data_in35;
  wire [7:0] data_in35;
  input [7:0] data_in36;
  wire [7:0] data_in36;
  input [7:0] data_in37;
  wire [7:0] data_in37;
  input [7:0] data_in38;
  wire [7:0] data_in38;
  input [7:0] data_in39;
  wire [7:0] data_in39;
  input [7:0] data_in40;
  wire [7:0] data_in40;
  input [7:0] data_in41;
  wire [7:0] data_in41;
  input [7:0] data_in42;
  wire [7:0] data_in42;
  input [7:0] data_in43;
  wire [7:0] data_in43;
  input [7:0] data_in44;
  wire [7:0] data_in44;
  input [7:0] data_in45;
  wire [7:0] data_in45;
  input [7:0] data_in46;
  wire [7:0] data_in46;
  input [7:0] data_in49;
  wire [7:0] data_in49;
  input [7:0] data_in50;
  wire [7:0] data_in50;
  input [7:0] data_in51;
  wire [7:0] data_in51;
  input [7:0] data_in52;
  wire [7:0] data_in52;
  input [7:0] data_in53;
  wire [7:0] data_in53;
  input [7:0] data_in54;
  wire [7:0] data_in54;
  input [7:0] data_in55;
  wire [7:0] data_in55;
  input [7:0] data_in56;
  wire [7:0] data_in56;
  input [7:0] data_in57;
  wire [7:0] data_in57;
  input [7:0] data_in58;
  wire [7:0] data_in58;
  input [7:0] data_in59;
  wire [7:0] data_in59;
  input [7:0] data_in60;
  wire [7:0] data_in60;
  input [7:0] data_in61;
  wire [7:0] data_in61;
  input [7:0] data_in62;
  wire [7:0] data_in62;
  input [7:0] data_in65;
  wire [7:0] data_in65;
  input [7:0] data_in66;
  wire [7:0] data_in66;
  input [7:0] data_in67;
  wire [7:0] data_in67;
  input [7:0] data_in68;
  wire [7:0] data_in68;
  input [7:0] data_in69;
  wire [7:0] data_in69;
  input [7:0] data_in70;
  wire [7:0] data_in70;
  input [7:0] data_in71;
  wire [7:0] data_in71;
  input [7:0] data_in72;
  wire [7:0] data_in72;
  input [7:0] data_in73;
  wire [7:0] data_in73;
  input [7:0] data_in74;
  wire [7:0] data_in74;
  input [7:0] data_in75;
  wire [7:0] data_in75;
  input [7:0] data_in76;
  wire [7:0] data_in76;
  input [7:0] data_in77;
  wire [7:0] data_in77;
  input [7:0] data_in78;
  wire [7:0] data_in78;
  input [7:0] data_in81;
  wire [7:0] data_in81;
  input [7:0] data_in82;
  wire [7:0] data_in82;
  input [7:0] data_in83;
  wire [7:0] data_in83;
  input [7:0] data_in84;
  wire [7:0] data_in84;
  input [7:0] data_in85;
  wire [7:0] data_in85;
  input [7:0] data_in86;
  wire [7:0] data_in86;
  input [7:0] data_in87;
  wire [7:0] data_in87;
  input [7:0] data_in88;
  wire [7:0] data_in88;
  input [7:0] data_in89;
  wire [7:0] data_in89;
  input [7:0] data_in90;
  wire [7:0] data_in90;
  input [7:0] data_in91;
  wire [7:0] data_in91;
  input [7:0] data_in92;
  wire [7:0] data_in92;
  input [7:0] data_in93;
  wire [7:0] data_in93;
  input [7:0] data_in94;
  wire [7:0] data_in94;
  input [7:0] data_in97;
  wire [7:0] data_in97;
  input [7:0] data_in98;
  wire [7:0] data_in98;
  input [7:0] data_in99;
  wire [7:0] data_in99;
  input [7:0] data_in100;
  wire [7:0] data_in100;
  input [7:0] data_in101;
  wire [7:0] data_in101;
  input [7:0] data_in102;
  wire [7:0] data_in102;
  input [7:0] data_in103;
  wire [7:0] data_in103;
  input [7:0] data_in104;
  wire [7:0] data_in104;
  input [7:0] data_in105;
  wire [7:0] data_in105;
  input [7:0] data_in106;
  wire [7:0] data_in106;
  input [7:0] data_in107;
  wire [7:0] data_in107;
  input [7:0] data_in108;
  wire [7:0] data_in108;
  input [7:0] data_in109;
  wire [7:0] data_in109;
  input [7:0] data_in110;
  wire [7:0] data_in110;
  output [7:0] data_out17;
  wire [7:0] data_out17;
  output [7:0] data_out18;
  wire [7:0] data_out18;
  output [7:0] data_out19;
  wire [7:0] data_out19;
  output [7:0] data_out20;
  wire [7:0] data_out20;
  output [7:0] data_out21;
  wire [7:0] data_out21;
  output [7:0] data_out22;
  wire [7:0] data_out22;
  output [7:0] data_out23;
  wire [7:0] data_out23;
  output [7:0] data_out24;
  wire [7:0] data_out24;
  output [7:0] data_out25;
  wire [7:0] data_out25;
  output [7:0] data_out26;
  wire [7:0] data_out26;
  output [7:0] data_out27;
  wire [7:0] data_out27;
  output [7:0] data_out28;
  wire [7:0] data_out28;
  output [7:0] data_out29;
  wire [7:0] data_out29;
  output [7:0] data_out30;
  wire [7:0] data_out30;
  output [7:0] data_out33;
  wire [7:0] data_out33;
  output [7:0] data_out34;
  wire [7:0] data_out34;
  output [7:0] data_out35;
  wire [7:0] data_out35;
  output [7:0] data_out36;
  wire [7:0] data_out36;
  output [7:0] data_out37;
  wire [7:0] data_out37;
  output [7:0] data_out38;
  wire [7:0] data_out38;
  output [7:0] data_out39;
  wire [7:0] data_out39;
  output [7:0] data_out40;
  wire [7:0] data_out40;
  output [7:0] data_out41;
  wire [7:0] data_out41;
  output [7:0] data_out42;
  wire [7:0] data_out42;
  output [7:0] data_out43;
  wire [7:0] data_out43;
  output [7:0] data_out44;
  wire [7:0] data_out44;
  output [7:0] data_out45;
  wire [7:0] data_out45;
  output [7:0] data_out46;
  wire [7:0] data_out46;
  output [7:0] data_out49;
  wire [7:0] data_out49;
  output [7:0] data_out50;
  wire [7:0] data_out50;
  output [7:0] data_out51;
  wire [7:0] data_out51;
  output [7:0] data_out52;
  wire [7:0] data_out52;
  output [7:0] data_out53;
  wire [7:0] data_out53;
  output [7:0] data_out54;
  wire [7:0] data_out54;
  output [7:0] data_out55;
  wire [7:0] data_out55;
  output [7:0] data_out56;
  wire [7:0] data_out56;
  output [7:0] data_out57;
  wire [7:0] data_out57;
  output [7:0] data_out58;
  wire [7:0] data_out58;
  output [7:0] data_out59;
  wire [7:0] data_out59;
  output [7:0] data_out60;
  wire [7:0] data_out60;
  output [7:0] data_out61;
  wire [7:0] data_out61;
  output [7:0] data_out62;
  wire [7:0] data_out62;
  output [7:0] data_out65;
  wire [7:0] data_out65;
  output [7:0] data_out66;
  wire [7:0] data_out66;
  output [7:0] data_out67;
  wire [7:0] data_out67;
  output [7:0] data_out68;
  wire [7:0] data_out68;
  output [7:0] data_out69;
  wire [7:0] data_out69;
  output [7:0] data_out70;
  wire [7:0] data_out70;
  output [7:0] data_out71;
  wire [7:0] data_out71;
  output [7:0] data_out72;
  wire [7:0] data_out72;
  output [7:0] data_out73;
  wire [7:0] data_out73;
  output [7:0] data_out74;
  wire [7:0] data_out74;
  output [7:0] data_out75;
  wire [7:0] data_out75;
  output [7:0] data_out76;
  wire [7:0] data_out76;
  output [7:0] data_out77;
  wire [7:0] data_out77;
  output [7:0] data_out78;
  wire [7:0] data_out78;
  output [7:0] data_out81;
  wire [7:0] data_out81;
  output [7:0] data_out82;
  wire [7:0] data_out82;
  output [7:0] data_out83;
  wire [7:0] data_out83;
  output [7:0] data_out84;
  wire [7:0] data_out84;
  output [7:0] data_out85;
  wire [7:0] data_out85;
  output [7:0] data_out86;
  wire [7:0] data_out86;
  output [7:0] data_out87;
  wire [7:0] data_out87;
  output [7:0] data_out88;
  wire [7:0] data_out88;
  output [7:0] data_out89;
  wire [7:0] data_out89;
  output [7:0] data_out90;
  wire [7:0] data_out90;
  output [7:0] data_out91;
  wire [7:0] data_out91;
  output [7:0] data_out92;
  wire [7:0] data_out92;
  output [7:0] data_out93;
  wire [7:0] data_out93;
  output [7:0] data_out94;
  wire [7:0] data_out94;
  output [7:0] data_out97;
  wire [7:0] data_out97;
  output [7:0] data_out98;
  wire [7:0] data_out98;
  output [7:0] data_out99;
  wire [7:0] data_out99;
  output [7:0] data_out100;
  wire [7:0] data_out100;
  output [7:0] data_out101;
  wire [7:0] data_out101;
  output [7:0] data_out102;
  wire [7:0] data_out102;
  output [7:0] data_out103;
  wire [7:0] data_out103;
  output [7:0] data_out104;
  wire [7:0] data_out104;
  output [7:0] data_out105;
  wire [7:0] data_out105;
  output [7:0] data_out106;
  wire [7:0] data_out106;
  output [7:0] data_out107;
  wire [7:0] data_out107;
  output [7:0] data_out108;
  wire [7:0] data_out108;
  output [7:0] data_out109;
  wire [7:0] data_out109;
  output [7:0] data_out110;
  wire [7:0] data_out110;
  output [7:0] startplot;
  wire [7:0] startplot;
  output [7:0] goalplot;
  wire [7:0] goalplot;
  input in_do;
  wire in_do;
  output out_do;
  wire out_do;
  output out_data;
  wire out_data;
  reg [7:0] startplot_reg;
  reg [7:0] goalplot_reg;
  wire [7:0] startplot_wire;
  wire [7:0] goalplot_wire;
  wire [7:0] _seach_blockx_map_block;
  wire [7:0] _seach_blockx_now;
  wire [7:0] _seach_blockx_start;
  wire [7:0] _seach_blockx_goal;
  wire [7:0] _seach_blockx_data_out;
  wire _seach_blockx_in_do;
  wire _seach_blockx_p_reset;
  wire _seach_blockx_m_clock;
  wire [7:0] _seach_blockx_195_map_block;
  wire [7:0] _seach_blockx_195_now;
  wire [7:0] _seach_blockx_195_start;
  wire [7:0] _seach_blockx_195_goal;
  wire [7:0] _seach_blockx_195_data_out;
  wire _seach_blockx_195_in_do;
  wire _seach_blockx_195_p_reset;
  wire _seach_blockx_195_m_clock;
  wire [7:0] _seach_blockx_194_map_block;
  wire [7:0] _seach_blockx_194_now;
  wire [7:0] _seach_blockx_194_start;
  wire [7:0] _seach_blockx_194_goal;
  wire [7:0] _seach_blockx_194_data_out;
  wire _seach_blockx_194_in_do;
  wire _seach_blockx_194_p_reset;
  wire _seach_blockx_194_m_clock;
  wire [7:0] _seach_blockx_193_map_block;
  wire [7:0] _seach_blockx_193_now;
  wire [7:0] _seach_blockx_193_start;
  wire [7:0] _seach_blockx_193_goal;
  wire [7:0] _seach_blockx_193_data_out;
  wire _seach_blockx_193_in_do;
  wire _seach_blockx_193_p_reset;
  wire _seach_blockx_193_m_clock;
  wire [7:0] _seach_blockx_192_map_block;
  wire [7:0] _seach_blockx_192_now;
  wire [7:0] _seach_blockx_192_start;
  wire [7:0] _seach_blockx_192_goal;
  wire [7:0] _seach_blockx_192_data_out;
  wire _seach_blockx_192_in_do;
  wire _seach_blockx_192_p_reset;
  wire _seach_blockx_192_m_clock;
  wire [7:0] _seach_blockx_191_map_block;
  wire [7:0] _seach_blockx_191_now;
  wire [7:0] _seach_blockx_191_start;
  wire [7:0] _seach_blockx_191_goal;
  wire [7:0] _seach_blockx_191_data_out;
  wire _seach_blockx_191_in_do;
  wire _seach_blockx_191_p_reset;
  wire _seach_blockx_191_m_clock;
  wire [7:0] _seach_blockx_190_map_block;
  wire [7:0] _seach_blockx_190_now;
  wire [7:0] _seach_blockx_190_start;
  wire [7:0] _seach_blockx_190_goal;
  wire [7:0] _seach_blockx_190_data_out;
  wire _seach_blockx_190_in_do;
  wire _seach_blockx_190_p_reset;
  wire _seach_blockx_190_m_clock;
  wire [7:0] _seach_blockx_189_map_block;
  wire [7:0] _seach_blockx_189_now;
  wire [7:0] _seach_blockx_189_start;
  wire [7:0] _seach_blockx_189_goal;
  wire [7:0] _seach_blockx_189_data_out;
  wire _seach_blockx_189_in_do;
  wire _seach_blockx_189_p_reset;
  wire _seach_blockx_189_m_clock;
  wire [7:0] _seach_blockx_188_map_block;
  wire [7:0] _seach_blockx_188_now;
  wire [7:0] _seach_blockx_188_start;
  wire [7:0] _seach_blockx_188_goal;
  wire [7:0] _seach_blockx_188_data_out;
  wire _seach_blockx_188_in_do;
  wire _seach_blockx_188_p_reset;
  wire _seach_blockx_188_m_clock;
  wire [7:0] _seach_blockx_187_map_block;
  wire [7:0] _seach_blockx_187_now;
  wire [7:0] _seach_blockx_187_start;
  wire [7:0] _seach_blockx_187_goal;
  wire [7:0] _seach_blockx_187_data_out;
  wire _seach_blockx_187_in_do;
  wire _seach_blockx_187_p_reset;
  wire _seach_blockx_187_m_clock;
  wire [7:0] _seach_blockx_186_map_block;
  wire [7:0] _seach_blockx_186_now;
  wire [7:0] _seach_blockx_186_start;
  wire [7:0] _seach_blockx_186_goal;
  wire [7:0] _seach_blockx_186_data_out;
  wire _seach_blockx_186_in_do;
  wire _seach_blockx_186_p_reset;
  wire _seach_blockx_186_m_clock;
  wire [7:0] _seach_blockx_185_map_block;
  wire [7:0] _seach_blockx_185_now;
  wire [7:0] _seach_blockx_185_start;
  wire [7:0] _seach_blockx_185_goal;
  wire [7:0] _seach_blockx_185_data_out;
  wire _seach_blockx_185_in_do;
  wire _seach_blockx_185_p_reset;
  wire _seach_blockx_185_m_clock;
  wire [7:0] _seach_blockx_184_map_block;
  wire [7:0] _seach_blockx_184_now;
  wire [7:0] _seach_blockx_184_start;
  wire [7:0] _seach_blockx_184_goal;
  wire [7:0] _seach_blockx_184_data_out;
  wire _seach_blockx_184_in_do;
  wire _seach_blockx_184_p_reset;
  wire _seach_blockx_184_m_clock;
  wire [7:0] _seach_blockx_183_map_block;
  wire [7:0] _seach_blockx_183_now;
  wire [7:0] _seach_blockx_183_start;
  wire [7:0] _seach_blockx_183_goal;
  wire [7:0] _seach_blockx_183_data_out;
  wire _seach_blockx_183_in_do;
  wire _seach_blockx_183_p_reset;
  wire _seach_blockx_183_m_clock;
  wire [7:0] _seach_blockx_182_map_block;
  wire [7:0] _seach_blockx_182_now;
  wire [7:0] _seach_blockx_182_start;
  wire [7:0] _seach_blockx_182_goal;
  wire [7:0] _seach_blockx_182_data_out;
  wire _seach_blockx_182_in_do;
  wire _seach_blockx_182_p_reset;
  wire _seach_blockx_182_m_clock;
  wire [7:0] _seach_blockx_181_map_block;
  wire [7:0] _seach_blockx_181_now;
  wire [7:0] _seach_blockx_181_start;
  wire [7:0] _seach_blockx_181_goal;
  wire [7:0] _seach_blockx_181_data_out;
  wire _seach_blockx_181_in_do;
  wire _seach_blockx_181_p_reset;
  wire _seach_blockx_181_m_clock;
  wire [7:0] _seach_blockx_180_map_block;
  wire [7:0] _seach_blockx_180_now;
  wire [7:0] _seach_blockx_180_start;
  wire [7:0] _seach_blockx_180_goal;
  wire [7:0] _seach_blockx_180_data_out;
  wire _seach_blockx_180_in_do;
  wire _seach_blockx_180_p_reset;
  wire _seach_blockx_180_m_clock;
  wire [7:0] _seach_blockx_179_map_block;
  wire [7:0] _seach_blockx_179_now;
  wire [7:0] _seach_blockx_179_start;
  wire [7:0] _seach_blockx_179_goal;
  wire [7:0] _seach_blockx_179_data_out;
  wire _seach_blockx_179_in_do;
  wire _seach_blockx_179_p_reset;
  wire _seach_blockx_179_m_clock;
  wire [7:0] _seach_blockx_178_map_block;
  wire [7:0] _seach_blockx_178_now;
  wire [7:0] _seach_blockx_178_start;
  wire [7:0] _seach_blockx_178_goal;
  wire [7:0] _seach_blockx_178_data_out;
  wire _seach_blockx_178_in_do;
  wire _seach_blockx_178_p_reset;
  wire _seach_blockx_178_m_clock;
  wire [7:0] _seach_blockx_177_map_block;
  wire [7:0] _seach_blockx_177_now;
  wire [7:0] _seach_blockx_177_start;
  wire [7:0] _seach_blockx_177_goal;
  wire [7:0] _seach_blockx_177_data_out;
  wire _seach_blockx_177_in_do;
  wire _seach_blockx_177_p_reset;
  wire _seach_blockx_177_m_clock;
  wire [7:0] _seach_blockx_176_map_block;
  wire [7:0] _seach_blockx_176_now;
  wire [7:0] _seach_blockx_176_start;
  wire [7:0] _seach_blockx_176_goal;
  wire [7:0] _seach_blockx_176_data_out;
  wire _seach_blockx_176_in_do;
  wire _seach_blockx_176_p_reset;
  wire _seach_blockx_176_m_clock;
  wire [7:0] _seach_blockx_175_map_block;
  wire [7:0] _seach_blockx_175_now;
  wire [7:0] _seach_blockx_175_start;
  wire [7:0] _seach_blockx_175_goal;
  wire [7:0] _seach_blockx_175_data_out;
  wire _seach_blockx_175_in_do;
  wire _seach_blockx_175_p_reset;
  wire _seach_blockx_175_m_clock;
  wire [7:0] _seach_blockx_174_map_block;
  wire [7:0] _seach_blockx_174_now;
  wire [7:0] _seach_blockx_174_start;
  wire [7:0] _seach_blockx_174_goal;
  wire [7:0] _seach_blockx_174_data_out;
  wire _seach_blockx_174_in_do;
  wire _seach_blockx_174_p_reset;
  wire _seach_blockx_174_m_clock;
  wire [7:0] _seach_blockx_173_map_block;
  wire [7:0] _seach_blockx_173_now;
  wire [7:0] _seach_blockx_173_start;
  wire [7:0] _seach_blockx_173_goal;
  wire [7:0] _seach_blockx_173_data_out;
  wire _seach_blockx_173_in_do;
  wire _seach_blockx_173_p_reset;
  wire _seach_blockx_173_m_clock;
  wire [7:0] _seach_blockx_172_map_block;
  wire [7:0] _seach_blockx_172_now;
  wire [7:0] _seach_blockx_172_start;
  wire [7:0] _seach_blockx_172_goal;
  wire [7:0] _seach_blockx_172_data_out;
  wire _seach_blockx_172_in_do;
  wire _seach_blockx_172_p_reset;
  wire _seach_blockx_172_m_clock;
  wire [7:0] _seach_blockx_171_map_block;
  wire [7:0] _seach_blockx_171_now;
  wire [7:0] _seach_blockx_171_start;
  wire [7:0] _seach_blockx_171_goal;
  wire [7:0] _seach_blockx_171_data_out;
  wire _seach_blockx_171_in_do;
  wire _seach_blockx_171_p_reset;
  wire _seach_blockx_171_m_clock;
  wire [7:0] _seach_blockx_170_map_block;
  wire [7:0] _seach_blockx_170_now;
  wire [7:0] _seach_blockx_170_start;
  wire [7:0] _seach_blockx_170_goal;
  wire [7:0] _seach_blockx_170_data_out;
  wire _seach_blockx_170_in_do;
  wire _seach_blockx_170_p_reset;
  wire _seach_blockx_170_m_clock;
  wire [7:0] _seach_blockx_169_map_block;
  wire [7:0] _seach_blockx_169_now;
  wire [7:0] _seach_blockx_169_start;
  wire [7:0] _seach_blockx_169_goal;
  wire [7:0] _seach_blockx_169_data_out;
  wire _seach_blockx_169_in_do;
  wire _seach_blockx_169_p_reset;
  wire _seach_blockx_169_m_clock;
  wire [7:0] _seach_blockx_168_map_block;
  wire [7:0] _seach_blockx_168_now;
  wire [7:0] _seach_blockx_168_start;
  wire [7:0] _seach_blockx_168_goal;
  wire [7:0] _seach_blockx_168_data_out;
  wire _seach_blockx_168_in_do;
  wire _seach_blockx_168_p_reset;
  wire _seach_blockx_168_m_clock;
  wire [7:0] _seach_blockx_167_map_block;
  wire [7:0] _seach_blockx_167_now;
  wire [7:0] _seach_blockx_167_start;
  wire [7:0] _seach_blockx_167_goal;
  wire [7:0] _seach_blockx_167_data_out;
  wire _seach_blockx_167_in_do;
  wire _seach_blockx_167_p_reset;
  wire _seach_blockx_167_m_clock;
  wire [7:0] _seach_blockx_166_map_block;
  wire [7:0] _seach_blockx_166_now;
  wire [7:0] _seach_blockx_166_start;
  wire [7:0] _seach_blockx_166_goal;
  wire [7:0] _seach_blockx_166_data_out;
  wire _seach_blockx_166_in_do;
  wire _seach_blockx_166_p_reset;
  wire _seach_blockx_166_m_clock;
  wire [7:0] _seach_blockx_165_map_block;
  wire [7:0] _seach_blockx_165_now;
  wire [7:0] _seach_blockx_165_start;
  wire [7:0] _seach_blockx_165_goal;
  wire [7:0] _seach_blockx_165_data_out;
  wire _seach_blockx_165_in_do;
  wire _seach_blockx_165_p_reset;
  wire _seach_blockx_165_m_clock;
  wire [7:0] _seach_blockx_164_map_block;
  wire [7:0] _seach_blockx_164_now;
  wire [7:0] _seach_blockx_164_start;
  wire [7:0] _seach_blockx_164_goal;
  wire [7:0] _seach_blockx_164_data_out;
  wire _seach_blockx_164_in_do;
  wire _seach_blockx_164_p_reset;
  wire _seach_blockx_164_m_clock;
  wire [7:0] _seach_blockx_163_map_block;
  wire [7:0] _seach_blockx_163_now;
  wire [7:0] _seach_blockx_163_start;
  wire [7:0] _seach_blockx_163_goal;
  wire [7:0] _seach_blockx_163_data_out;
  wire _seach_blockx_163_in_do;
  wire _seach_blockx_163_p_reset;
  wire _seach_blockx_163_m_clock;
  wire [7:0] _seach_blockx_162_map_block;
  wire [7:0] _seach_blockx_162_now;
  wire [7:0] _seach_blockx_162_start;
  wire [7:0] _seach_blockx_162_goal;
  wire [7:0] _seach_blockx_162_data_out;
  wire _seach_blockx_162_in_do;
  wire _seach_blockx_162_p_reset;
  wire _seach_blockx_162_m_clock;
  wire [7:0] _seach_blockx_161_map_block;
  wire [7:0] _seach_blockx_161_now;
  wire [7:0] _seach_blockx_161_start;
  wire [7:0] _seach_blockx_161_goal;
  wire [7:0] _seach_blockx_161_data_out;
  wire _seach_blockx_161_in_do;
  wire _seach_blockx_161_p_reset;
  wire _seach_blockx_161_m_clock;
  wire [7:0] _seach_blockx_160_map_block;
  wire [7:0] _seach_blockx_160_now;
  wire [7:0] _seach_blockx_160_start;
  wire [7:0] _seach_blockx_160_goal;
  wire [7:0] _seach_blockx_160_data_out;
  wire _seach_blockx_160_in_do;
  wire _seach_blockx_160_p_reset;
  wire _seach_blockx_160_m_clock;
  wire [7:0] _seach_blockx_159_map_block;
  wire [7:0] _seach_blockx_159_now;
  wire [7:0] _seach_blockx_159_start;
  wire [7:0] _seach_blockx_159_goal;
  wire [7:0] _seach_blockx_159_data_out;
  wire _seach_blockx_159_in_do;
  wire _seach_blockx_159_p_reset;
  wire _seach_blockx_159_m_clock;
  wire [7:0] _seach_blockx_158_map_block;
  wire [7:0] _seach_blockx_158_now;
  wire [7:0] _seach_blockx_158_start;
  wire [7:0] _seach_blockx_158_goal;
  wire [7:0] _seach_blockx_158_data_out;
  wire _seach_blockx_158_in_do;
  wire _seach_blockx_158_p_reset;
  wire _seach_blockx_158_m_clock;
  wire [7:0] _seach_blockx_157_map_block;
  wire [7:0] _seach_blockx_157_now;
  wire [7:0] _seach_blockx_157_start;
  wire [7:0] _seach_blockx_157_goal;
  wire [7:0] _seach_blockx_157_data_out;
  wire _seach_blockx_157_in_do;
  wire _seach_blockx_157_p_reset;
  wire _seach_blockx_157_m_clock;
  wire [7:0] _seach_blockx_156_map_block;
  wire [7:0] _seach_blockx_156_now;
  wire [7:0] _seach_blockx_156_start;
  wire [7:0] _seach_blockx_156_goal;
  wire [7:0] _seach_blockx_156_data_out;
  wire _seach_blockx_156_in_do;
  wire _seach_blockx_156_p_reset;
  wire _seach_blockx_156_m_clock;
  wire [7:0] _seach_blockx_155_map_block;
  wire [7:0] _seach_blockx_155_now;
  wire [7:0] _seach_blockx_155_start;
  wire [7:0] _seach_blockx_155_goal;
  wire [7:0] _seach_blockx_155_data_out;
  wire _seach_blockx_155_in_do;
  wire _seach_blockx_155_p_reset;
  wire _seach_blockx_155_m_clock;
  wire [7:0] _seach_blockx_154_map_block;
  wire [7:0] _seach_blockx_154_now;
  wire [7:0] _seach_blockx_154_start;
  wire [7:0] _seach_blockx_154_goal;
  wire [7:0] _seach_blockx_154_data_out;
  wire _seach_blockx_154_in_do;
  wire _seach_blockx_154_p_reset;
  wire _seach_blockx_154_m_clock;
  wire [7:0] _seach_blockx_153_map_block;
  wire [7:0] _seach_blockx_153_now;
  wire [7:0] _seach_blockx_153_start;
  wire [7:0] _seach_blockx_153_goal;
  wire [7:0] _seach_blockx_153_data_out;
  wire _seach_blockx_153_in_do;
  wire _seach_blockx_153_p_reset;
  wire _seach_blockx_153_m_clock;
  wire [7:0] _seach_blockx_152_map_block;
  wire [7:0] _seach_blockx_152_now;
  wire [7:0] _seach_blockx_152_start;
  wire [7:0] _seach_blockx_152_goal;
  wire [7:0] _seach_blockx_152_data_out;
  wire _seach_blockx_152_in_do;
  wire _seach_blockx_152_p_reset;
  wire _seach_blockx_152_m_clock;
  wire [7:0] _seach_blockx_151_map_block;
  wire [7:0] _seach_blockx_151_now;
  wire [7:0] _seach_blockx_151_start;
  wire [7:0] _seach_blockx_151_goal;
  wire [7:0] _seach_blockx_151_data_out;
  wire _seach_blockx_151_in_do;
  wire _seach_blockx_151_p_reset;
  wire _seach_blockx_151_m_clock;
  wire [7:0] _seach_blockx_150_map_block;
  wire [7:0] _seach_blockx_150_now;
  wire [7:0] _seach_blockx_150_start;
  wire [7:0] _seach_blockx_150_goal;
  wire [7:0] _seach_blockx_150_data_out;
  wire _seach_blockx_150_in_do;
  wire _seach_blockx_150_p_reset;
  wire _seach_blockx_150_m_clock;
  wire [7:0] _seach_blockx_149_map_block;
  wire [7:0] _seach_blockx_149_now;
  wire [7:0] _seach_blockx_149_start;
  wire [7:0] _seach_blockx_149_goal;
  wire [7:0] _seach_blockx_149_data_out;
  wire _seach_blockx_149_in_do;
  wire _seach_blockx_149_p_reset;
  wire _seach_blockx_149_m_clock;
  wire [7:0] _seach_blockx_148_map_block;
  wire [7:0] _seach_blockx_148_now;
  wire [7:0] _seach_blockx_148_start;
  wire [7:0] _seach_blockx_148_goal;
  wire [7:0] _seach_blockx_148_data_out;
  wire _seach_blockx_148_in_do;
  wire _seach_blockx_148_p_reset;
  wire _seach_blockx_148_m_clock;
  wire [7:0] _seach_blockx_147_map_block;
  wire [7:0] _seach_blockx_147_now;
  wire [7:0] _seach_blockx_147_start;
  wire [7:0] _seach_blockx_147_goal;
  wire [7:0] _seach_blockx_147_data_out;
  wire _seach_blockx_147_in_do;
  wire _seach_blockx_147_p_reset;
  wire _seach_blockx_147_m_clock;
  wire [7:0] _seach_blockx_146_map_block;
  wire [7:0] _seach_blockx_146_now;
  wire [7:0] _seach_blockx_146_start;
  wire [7:0] _seach_blockx_146_goal;
  wire [7:0] _seach_blockx_146_data_out;
  wire _seach_blockx_146_in_do;
  wire _seach_blockx_146_p_reset;
  wire _seach_blockx_146_m_clock;
  wire [7:0] _seach_blockx_145_map_block;
  wire [7:0] _seach_blockx_145_now;
  wire [7:0] _seach_blockx_145_start;
  wire [7:0] _seach_blockx_145_goal;
  wire [7:0] _seach_blockx_145_data_out;
  wire _seach_blockx_145_in_do;
  wire _seach_blockx_145_p_reset;
  wire _seach_blockx_145_m_clock;
  wire [7:0] _seach_blockx_144_map_block;
  wire [7:0] _seach_blockx_144_now;
  wire [7:0] _seach_blockx_144_start;
  wire [7:0] _seach_blockx_144_goal;
  wire [7:0] _seach_blockx_144_data_out;
  wire _seach_blockx_144_in_do;
  wire _seach_blockx_144_p_reset;
  wire _seach_blockx_144_m_clock;
  wire [7:0] _seach_blockx_143_map_block;
  wire [7:0] _seach_blockx_143_now;
  wire [7:0] _seach_blockx_143_start;
  wire [7:0] _seach_blockx_143_goal;
  wire [7:0] _seach_blockx_143_data_out;
  wire _seach_blockx_143_in_do;
  wire _seach_blockx_143_p_reset;
  wire _seach_blockx_143_m_clock;
  wire [7:0] _seach_blockx_142_map_block;
  wire [7:0] _seach_blockx_142_now;
  wire [7:0] _seach_blockx_142_start;
  wire [7:0] _seach_blockx_142_goal;
  wire [7:0] _seach_blockx_142_data_out;
  wire _seach_blockx_142_in_do;
  wire _seach_blockx_142_p_reset;
  wire _seach_blockx_142_m_clock;
  wire [7:0] _seach_blockx_141_map_block;
  wire [7:0] _seach_blockx_141_now;
  wire [7:0] _seach_blockx_141_start;
  wire [7:0] _seach_blockx_141_goal;
  wire [7:0] _seach_blockx_141_data_out;
  wire _seach_blockx_141_in_do;
  wire _seach_blockx_141_p_reset;
  wire _seach_blockx_141_m_clock;
  wire [7:0] _seach_blockx_140_map_block;
  wire [7:0] _seach_blockx_140_now;
  wire [7:0] _seach_blockx_140_start;
  wire [7:0] _seach_blockx_140_goal;
  wire [7:0] _seach_blockx_140_data_out;
  wire _seach_blockx_140_in_do;
  wire _seach_blockx_140_p_reset;
  wire _seach_blockx_140_m_clock;
  wire [7:0] _seach_blockx_139_map_block;
  wire [7:0] _seach_blockx_139_now;
  wire [7:0] _seach_blockx_139_start;
  wire [7:0] _seach_blockx_139_goal;
  wire [7:0] _seach_blockx_139_data_out;
  wire _seach_blockx_139_in_do;
  wire _seach_blockx_139_p_reset;
  wire _seach_blockx_139_m_clock;
  wire [7:0] _seach_blockx_138_map_block;
  wire [7:0] _seach_blockx_138_now;
  wire [7:0] _seach_blockx_138_start;
  wire [7:0] _seach_blockx_138_goal;
  wire [7:0] _seach_blockx_138_data_out;
  wire _seach_blockx_138_in_do;
  wire _seach_blockx_138_p_reset;
  wire _seach_blockx_138_m_clock;
  wire [7:0] _seach_blockx_137_map_block;
  wire [7:0] _seach_blockx_137_now;
  wire [7:0] _seach_blockx_137_start;
  wire [7:0] _seach_blockx_137_goal;
  wire [7:0] _seach_blockx_137_data_out;
  wire _seach_blockx_137_in_do;
  wire _seach_blockx_137_p_reset;
  wire _seach_blockx_137_m_clock;
  wire [7:0] _seach_blockx_136_map_block;
  wire [7:0] _seach_blockx_136_now;
  wire [7:0] _seach_blockx_136_start;
  wire [7:0] _seach_blockx_136_goal;
  wire [7:0] _seach_blockx_136_data_out;
  wire _seach_blockx_136_in_do;
  wire _seach_blockx_136_p_reset;
  wire _seach_blockx_136_m_clock;
  wire [7:0] _seach_blockx_135_map_block;
  wire [7:0] _seach_blockx_135_now;
  wire [7:0] _seach_blockx_135_start;
  wire [7:0] _seach_blockx_135_goal;
  wire [7:0] _seach_blockx_135_data_out;
  wire _seach_blockx_135_in_do;
  wire _seach_blockx_135_p_reset;
  wire _seach_blockx_135_m_clock;
  wire [7:0] _seach_blockx_134_map_block;
  wire [7:0] _seach_blockx_134_now;
  wire [7:0] _seach_blockx_134_start;
  wire [7:0] _seach_blockx_134_goal;
  wire [7:0] _seach_blockx_134_data_out;
  wire _seach_blockx_134_in_do;
  wire _seach_blockx_134_p_reset;
  wire _seach_blockx_134_m_clock;
  wire [7:0] _seach_blockx_133_map_block;
  wire [7:0] _seach_blockx_133_now;
  wire [7:0] _seach_blockx_133_start;
  wire [7:0] _seach_blockx_133_goal;
  wire [7:0] _seach_blockx_133_data_out;
  wire _seach_blockx_133_in_do;
  wire _seach_blockx_133_p_reset;
  wire _seach_blockx_133_m_clock;
  wire [7:0] _seach_blockx_132_map_block;
  wire [7:0] _seach_blockx_132_now;
  wire [7:0] _seach_blockx_132_start;
  wire [7:0] _seach_blockx_132_goal;
  wire [7:0] _seach_blockx_132_data_out;
  wire _seach_blockx_132_in_do;
  wire _seach_blockx_132_p_reset;
  wire _seach_blockx_132_m_clock;
  wire [7:0] _seach_blockx_131_map_block;
  wire [7:0] _seach_blockx_131_now;
  wire [7:0] _seach_blockx_131_start;
  wire [7:0] _seach_blockx_131_goal;
  wire [7:0] _seach_blockx_131_data_out;
  wire _seach_blockx_131_in_do;
  wire _seach_blockx_131_p_reset;
  wire _seach_blockx_131_m_clock;
  wire [7:0] _seach_blockx_130_map_block;
  wire [7:0] _seach_blockx_130_now;
  wire [7:0] _seach_blockx_130_start;
  wire [7:0] _seach_blockx_130_goal;
  wire [7:0] _seach_blockx_130_data_out;
  wire _seach_blockx_130_in_do;
  wire _seach_blockx_130_p_reset;
  wire _seach_blockx_130_m_clock;
  wire [7:0] _seach_blockx_129_map_block;
  wire [7:0] _seach_blockx_129_now;
  wire [7:0] _seach_blockx_129_start;
  wire [7:0] _seach_blockx_129_goal;
  wire [7:0] _seach_blockx_129_data_out;
  wire _seach_blockx_129_in_do;
  wire _seach_blockx_129_p_reset;
  wire _seach_blockx_129_m_clock;
  wire [7:0] _seach_blockx_128_map_block;
  wire [7:0] _seach_blockx_128_now;
  wire [7:0] _seach_blockx_128_start;
  wire [7:0] _seach_blockx_128_goal;
  wire [7:0] _seach_blockx_128_data_out;
  wire _seach_blockx_128_in_do;
  wire _seach_blockx_128_p_reset;
  wire _seach_blockx_128_m_clock;
  wire [7:0] _seach_blockx_127_map_block;
  wire [7:0] _seach_blockx_127_now;
  wire [7:0] _seach_blockx_127_start;
  wire [7:0] _seach_blockx_127_goal;
  wire [7:0] _seach_blockx_127_data_out;
  wire _seach_blockx_127_in_do;
  wire _seach_blockx_127_p_reset;
  wire _seach_blockx_127_m_clock;
  wire [7:0] _seach_blockx_126_map_block;
  wire [7:0] _seach_blockx_126_now;
  wire [7:0] _seach_blockx_126_start;
  wire [7:0] _seach_blockx_126_goal;
  wire [7:0] _seach_blockx_126_data_out;
  wire _seach_blockx_126_in_do;
  wire _seach_blockx_126_p_reset;
  wire _seach_blockx_126_m_clock;
  wire [7:0] _seach_blockx_125_map_block;
  wire [7:0] _seach_blockx_125_now;
  wire [7:0] _seach_blockx_125_start;
  wire [7:0] _seach_blockx_125_goal;
  wire [7:0] _seach_blockx_125_data_out;
  wire _seach_blockx_125_in_do;
  wire _seach_blockx_125_p_reset;
  wire _seach_blockx_125_m_clock;
  wire [7:0] _seach_blockx_124_map_block;
  wire [7:0] _seach_blockx_124_now;
  wire [7:0] _seach_blockx_124_start;
  wire [7:0] _seach_blockx_124_goal;
  wire [7:0] _seach_blockx_124_data_out;
  wire _seach_blockx_124_in_do;
  wire _seach_blockx_124_p_reset;
  wire _seach_blockx_124_m_clock;
  wire [7:0] _seach_blockx_123_map_block;
  wire [7:0] _seach_blockx_123_now;
  wire [7:0] _seach_blockx_123_start;
  wire [7:0] _seach_blockx_123_goal;
  wire [7:0] _seach_blockx_123_data_out;
  wire _seach_blockx_123_in_do;
  wire _seach_blockx_123_p_reset;
  wire _seach_blockx_123_m_clock;
  wire [7:0] _seach_blockx_122_map_block;
  wire [7:0] _seach_blockx_122_now;
  wire [7:0] _seach_blockx_122_start;
  wire [7:0] _seach_blockx_122_goal;
  wire [7:0] _seach_blockx_122_data_out;
  wire _seach_blockx_122_in_do;
  wire _seach_blockx_122_p_reset;
  wire _seach_blockx_122_m_clock;
  wire [7:0] _seach_blockx_121_map_block;
  wire [7:0] _seach_blockx_121_now;
  wire [7:0] _seach_blockx_121_start;
  wire [7:0] _seach_blockx_121_goal;
  wire [7:0] _seach_blockx_121_data_out;
  wire _seach_blockx_121_in_do;
  wire _seach_blockx_121_p_reset;
  wire _seach_blockx_121_m_clock;
  wire [7:0] _seach_blockx_120_map_block;
  wire [7:0] _seach_blockx_120_now;
  wire [7:0] _seach_blockx_120_start;
  wire [7:0] _seach_blockx_120_goal;
  wire [7:0] _seach_blockx_120_data_out;
  wire _seach_blockx_120_in_do;
  wire _seach_blockx_120_p_reset;
  wire _seach_blockx_120_m_clock;
  wire [7:0] _seach_blockx_119_map_block;
  wire [7:0] _seach_blockx_119_now;
  wire [7:0] _seach_blockx_119_start;
  wire [7:0] _seach_blockx_119_goal;
  wire [7:0] _seach_blockx_119_data_out;
  wire _seach_blockx_119_in_do;
  wire _seach_blockx_119_p_reset;
  wire _seach_blockx_119_m_clock;
  wire [7:0] _seach_blockx_118_map_block;
  wire [7:0] _seach_blockx_118_now;
  wire [7:0] _seach_blockx_118_start;
  wire [7:0] _seach_blockx_118_goal;
  wire [7:0] _seach_blockx_118_data_out;
  wire _seach_blockx_118_in_do;
  wire _seach_blockx_118_p_reset;
  wire _seach_blockx_118_m_clock;
  wire [7:0] _seach_blockx_117_map_block;
  wire [7:0] _seach_blockx_117_now;
  wire [7:0] _seach_blockx_117_start;
  wire [7:0] _seach_blockx_117_goal;
  wire [7:0] _seach_blockx_117_data_out;
  wire _seach_blockx_117_in_do;
  wire _seach_blockx_117_p_reset;
  wire _seach_blockx_117_m_clock;
  wire [7:0] _seach_blockx_116_map_block;
  wire [7:0] _seach_blockx_116_now;
  wire [7:0] _seach_blockx_116_start;
  wire [7:0] _seach_blockx_116_goal;
  wire [7:0] _seach_blockx_116_data_out;
  wire _seach_blockx_116_in_do;
  wire _seach_blockx_116_p_reset;
  wire _seach_blockx_116_m_clock;
  wire [7:0] _seach_blockx_115_map_block;
  wire [7:0] _seach_blockx_115_now;
  wire [7:0] _seach_blockx_115_start;
  wire [7:0] _seach_blockx_115_goal;
  wire [7:0] _seach_blockx_115_data_out;
  wire _seach_blockx_115_in_do;
  wire _seach_blockx_115_p_reset;
  wire _seach_blockx_115_m_clock;
  wire [7:0] _seach_blockx_114_map_block;
  wire [7:0] _seach_blockx_114_now;
  wire [7:0] _seach_blockx_114_start;
  wire [7:0] _seach_blockx_114_goal;
  wire [7:0] _seach_blockx_114_data_out;
  wire _seach_blockx_114_in_do;
  wire _seach_blockx_114_p_reset;
  wire _seach_blockx_114_m_clock;
  wire [7:0] _seach_blockx_113_map_block;
  wire [7:0] _seach_blockx_113_now;
  wire [7:0] _seach_blockx_113_start;
  wire [7:0] _seach_blockx_113_goal;
  wire [7:0] _seach_blockx_113_data_out;
  wire _seach_blockx_113_in_do;
  wire _seach_blockx_113_p_reset;
  wire _seach_blockx_113_m_clock;
  wire [7:0] _seach_blockx_112_map_block;
  wire [7:0] _seach_blockx_112_now;
  wire [7:0] _seach_blockx_112_start;
  wire [7:0] _seach_blockx_112_goal;
  wire [7:0] _seach_blockx_112_data_out;
  wire _seach_blockx_112_in_do;
  wire _seach_blockx_112_p_reset;
  wire _seach_blockx_112_m_clock;
  wire [7:0] _seach_blockx_111_map_block;
  wire [7:0] _seach_blockx_111_now;
  wire [7:0] _seach_blockx_111_start;
  wire [7:0] _seach_blockx_111_goal;
  wire [7:0] _seach_blockx_111_data_out;
  wire _seach_blockx_111_in_do;
  wire _seach_blockx_111_p_reset;
  wire _seach_blockx_111_m_clock;
  wire [7:0] _seach_blockx_110_map_block;
  wire [7:0] _seach_blockx_110_now;
  wire [7:0] _seach_blockx_110_start;
  wire [7:0] _seach_blockx_110_goal;
  wire [7:0] _seach_blockx_110_data_out;
  wire _seach_blockx_110_in_do;
  wire _seach_blockx_110_p_reset;
  wire _seach_blockx_110_m_clock;
  wire [7:0] _seach_blockx_109_map_block;
  wire [7:0] _seach_blockx_109_now;
  wire [7:0] _seach_blockx_109_start;
  wire [7:0] _seach_blockx_109_goal;
  wire [7:0] _seach_blockx_109_data_out;
  wire _seach_blockx_109_in_do;
  wire _seach_blockx_109_p_reset;
  wire _seach_blockx_109_m_clock;
  wire [7:0] _seach_blockx_108_map_block;
  wire [7:0] _seach_blockx_108_now;
  wire [7:0] _seach_blockx_108_start;
  wire [7:0] _seach_blockx_108_goal;
  wire [7:0] _seach_blockx_108_data_out;
  wire _seach_blockx_108_in_do;
  wire _seach_blockx_108_p_reset;
  wire _seach_blockx_108_m_clock;
  wire [7:0] _seach_blockx_107_map_block;
  wire [7:0] _seach_blockx_107_now;
  wire [7:0] _seach_blockx_107_start;
  wire [7:0] _seach_blockx_107_goal;
  wire [7:0] _seach_blockx_107_data_out;
  wire _seach_blockx_107_in_do;
  wire _seach_blockx_107_p_reset;
  wire _seach_blockx_107_m_clock;
  wire [7:0] _seach_blockx_106_map_block;
  wire [7:0] _seach_blockx_106_now;
  wire [7:0] _seach_blockx_106_start;
  wire [7:0] _seach_blockx_106_goal;
  wire [7:0] _seach_blockx_106_data_out;
  wire _seach_blockx_106_in_do;
  wire _seach_blockx_106_p_reset;
  wire _seach_blockx_106_m_clock;
  wire [7:0] _seach_blockx_105_map_block;
  wire [7:0] _seach_blockx_105_now;
  wire [7:0] _seach_blockx_105_start;
  wire [7:0] _seach_blockx_105_goal;
  wire [7:0] _seach_blockx_105_data_out;
  wire _seach_blockx_105_in_do;
  wire _seach_blockx_105_p_reset;
  wire _seach_blockx_105_m_clock;
  wire [7:0] _seach_blockx_104_map_block;
  wire [7:0] _seach_blockx_104_now;
  wire [7:0] _seach_blockx_104_start;
  wire [7:0] _seach_blockx_104_goal;
  wire [7:0] _seach_blockx_104_data_out;
  wire _seach_blockx_104_in_do;
  wire _seach_blockx_104_p_reset;
  wire _seach_blockx_104_m_clock;
  wire [7:0] _seach_blockx_103_map_block;
  wire [7:0] _seach_blockx_103_now;
  wire [7:0] _seach_blockx_103_start;
  wire [7:0] _seach_blockx_103_goal;
  wire [7:0] _seach_blockx_103_data_out;
  wire _seach_blockx_103_in_do;
  wire _seach_blockx_103_p_reset;
  wire _seach_blockx_103_m_clock;
  wire [7:0] _seach_blockx_102_map_block;
  wire [7:0] _seach_blockx_102_now;
  wire [7:0] _seach_blockx_102_start;
  wire [7:0] _seach_blockx_102_goal;
  wire [7:0] _seach_blockx_102_data_out;
  wire _seach_blockx_102_in_do;
  wire _seach_blockx_102_p_reset;
  wire _seach_blockx_102_m_clock;
  wire [7:0] _seach_blockx_101_map_block;
  wire [7:0] _seach_blockx_101_now;
  wire [7:0] _seach_blockx_101_start;
  wire [7:0] _seach_blockx_101_goal;
  wire [7:0] _seach_blockx_101_data_out;
  wire _seach_blockx_101_in_do;
  wire _seach_blockx_101_p_reset;
  wire _seach_blockx_101_m_clock;
  wire [7:0] _seach_blockx_100_map_block;
  wire [7:0] _seach_blockx_100_now;
  wire [7:0] _seach_blockx_100_start;
  wire [7:0] _seach_blockx_100_goal;
  wire [7:0] _seach_blockx_100_data_out;
  wire _seach_blockx_100_in_do;
  wire _seach_blockx_100_p_reset;
  wire _seach_blockx_100_m_clock;
  wire [7:0] _seach_blockx_99_map_block;
  wire [7:0] _seach_blockx_99_now;
  wire [7:0] _seach_blockx_99_start;
  wire [7:0] _seach_blockx_99_goal;
  wire [7:0] _seach_blockx_99_data_out;
  wire _seach_blockx_99_in_do;
  wire _seach_blockx_99_p_reset;
  wire _seach_blockx_99_m_clock;
  wire [7:0] _seach_blockx_98_map_block;
  wire [7:0] _seach_blockx_98_now;
  wire [7:0] _seach_blockx_98_start;
  wire [7:0] _seach_blockx_98_goal;
  wire [7:0] _seach_blockx_98_data_out;
  wire _seach_blockx_98_in_do;
  wire _seach_blockx_98_p_reset;
  wire _seach_blockx_98_m_clock;
  wire [7:0] _seach_blockx_97_map_block;
  wire [7:0] _seach_blockx_97_now;
  wire [7:0] _seach_blockx_97_start;
  wire [7:0] _seach_blockx_97_goal;
  wire [7:0] _seach_blockx_97_data_out;
  wire _seach_blockx_97_in_do;
  wire _seach_blockx_97_p_reset;
  wire _seach_blockx_97_m_clock;
  wire [7:0] _seach_blockx_96_map_block;
  wire [7:0] _seach_blockx_96_now;
  wire [7:0] _seach_blockx_96_start;
  wire [7:0] _seach_blockx_96_goal;
  wire [7:0] _seach_blockx_96_data_out;
  wire _seach_blockx_96_in_do;
  wire _seach_blockx_96_p_reset;
  wire _seach_blockx_96_m_clock;
  wire [7:0] _seach_blockx_95_map_block;
  wire [7:0] _seach_blockx_95_now;
  wire [7:0] _seach_blockx_95_start;
  wire [7:0] _seach_blockx_95_goal;
  wire [7:0] _seach_blockx_95_data_out;
  wire _seach_blockx_95_in_do;
  wire _seach_blockx_95_p_reset;
  wire _seach_blockx_95_m_clock;
  wire [7:0] _seach_blockx_94_map_block;
  wire [7:0] _seach_blockx_94_now;
  wire [7:0] _seach_blockx_94_start;
  wire [7:0] _seach_blockx_94_goal;
  wire [7:0] _seach_blockx_94_data_out;
  wire _seach_blockx_94_in_do;
  wire _seach_blockx_94_p_reset;
  wire _seach_blockx_94_m_clock;
  wire [7:0] _seach_blockx_93_map_block;
  wire [7:0] _seach_blockx_93_now;
  wire [7:0] _seach_blockx_93_start;
  wire [7:0] _seach_blockx_93_goal;
  wire [7:0] _seach_blockx_93_data_out;
  wire _seach_blockx_93_in_do;
  wire _seach_blockx_93_p_reset;
  wire _seach_blockx_93_m_clock;
  wire [7:0] _seach_blockx_92_map_block;
  wire [7:0] _seach_blockx_92_now;
  wire [7:0] _seach_blockx_92_start;
  wire [7:0] _seach_blockx_92_goal;
  wire [7:0] _seach_blockx_92_data_out;
  wire _seach_blockx_92_in_do;
  wire _seach_blockx_92_p_reset;
  wire _seach_blockx_92_m_clock;
  wire [7:0] _seach_blockx_91_map_block;
  wire [7:0] _seach_blockx_91_now;
  wire [7:0] _seach_blockx_91_start;
  wire [7:0] _seach_blockx_91_goal;
  wire [7:0] _seach_blockx_91_data_out;
  wire _seach_blockx_91_in_do;
  wire _seach_blockx_91_p_reset;
  wire _seach_blockx_91_m_clock;
  wire [7:0] _seach_blockx_90_map_block;
  wire [7:0] _seach_blockx_90_now;
  wire [7:0] _seach_blockx_90_start;
  wire [7:0] _seach_blockx_90_goal;
  wire [7:0] _seach_blockx_90_data_out;
  wire _seach_blockx_90_in_do;
  wire _seach_blockx_90_p_reset;
  wire _seach_blockx_90_m_clock;
  wire [7:0] _seach_blockx_89_map_block;
  wire [7:0] _seach_blockx_89_now;
  wire [7:0] _seach_blockx_89_start;
  wire [7:0] _seach_blockx_89_goal;
  wire [7:0] _seach_blockx_89_data_out;
  wire _seach_blockx_89_in_do;
  wire _seach_blockx_89_p_reset;
  wire _seach_blockx_89_m_clock;
  wire [7:0] _seach_blockx_88_map_block;
  wire [7:0] _seach_blockx_88_now;
  wire [7:0] _seach_blockx_88_start;
  wire [7:0] _seach_blockx_88_goal;
  wire [7:0] _seach_blockx_88_data_out;
  wire _seach_blockx_88_in_do;
  wire _seach_blockx_88_p_reset;
  wire _seach_blockx_88_m_clock;
  wire [7:0] _seach_blockx_87_map_block;
  wire [7:0] _seach_blockx_87_now;
  wire [7:0] _seach_blockx_87_start;
  wire [7:0] _seach_blockx_87_goal;
  wire [7:0] _seach_blockx_87_data_out;
  wire _seach_blockx_87_in_do;
  wire _seach_blockx_87_p_reset;
  wire _seach_blockx_87_m_clock;
  wire [7:0] _seach_blockx_86_map_block;
  wire [7:0] _seach_blockx_86_now;
  wire [7:0] _seach_blockx_86_start;
  wire [7:0] _seach_blockx_86_goal;
  wire [7:0] _seach_blockx_86_data_out;
  wire _seach_blockx_86_in_do;
  wire _seach_blockx_86_p_reset;
  wire _seach_blockx_86_m_clock;
  wire [7:0] _seach_blockx_85_map_block;
  wire [7:0] _seach_blockx_85_now;
  wire [7:0] _seach_blockx_85_start;
  wire [7:0] _seach_blockx_85_goal;
  wire [7:0] _seach_blockx_85_data_out;
  wire _seach_blockx_85_in_do;
  wire _seach_blockx_85_p_reset;
  wire _seach_blockx_85_m_clock;
  wire [7:0] _seach_blockx_84_map_block;
  wire [7:0] _seach_blockx_84_now;
  wire [7:0] _seach_blockx_84_start;
  wire [7:0] _seach_blockx_84_goal;
  wire [7:0] _seach_blockx_84_data_out;
  wire _seach_blockx_84_in_do;
  wire _seach_blockx_84_p_reset;
  wire _seach_blockx_84_m_clock;
  wire [7:0] _seach_blockx_83_map_block;
  wire [7:0] _seach_blockx_83_now;
  wire [7:0] _seach_blockx_83_start;
  wire [7:0] _seach_blockx_83_goal;
  wire [7:0] _seach_blockx_83_data_out;
  wire _seach_blockx_83_in_do;
  wire _seach_blockx_83_p_reset;
  wire _seach_blockx_83_m_clock;
  wire [7:0] _seach_blockx_82_map_block;
  wire [7:0] _seach_blockx_82_now;
  wire [7:0] _seach_blockx_82_start;
  wire [7:0] _seach_blockx_82_goal;
  wire [7:0] _seach_blockx_82_data_out;
  wire _seach_blockx_82_in_do;
  wire _seach_blockx_82_p_reset;
  wire _seach_blockx_82_m_clock;
  wire [7:0] _seach_blockx_81_map_block;
  wire [7:0] _seach_blockx_81_now;
  wire [7:0] _seach_blockx_81_start;
  wire [7:0] _seach_blockx_81_goal;
  wire [7:0] _seach_blockx_81_data_out;
  wire _seach_blockx_81_in_do;
  wire _seach_blockx_81_p_reset;
  wire _seach_blockx_81_m_clock;
  wire [7:0] _seach_blockx_80_map_block;
  wire [7:0] _seach_blockx_80_now;
  wire [7:0] _seach_blockx_80_start;
  wire [7:0] _seach_blockx_80_goal;
  wire [7:0] _seach_blockx_80_data_out;
  wire _seach_blockx_80_in_do;
  wire _seach_blockx_80_p_reset;
  wire _seach_blockx_80_m_clock;
  wire [7:0] _seach_blockx_79_map_block;
  wire [7:0] _seach_blockx_79_now;
  wire [7:0] _seach_blockx_79_start;
  wire [7:0] _seach_blockx_79_goal;
  wire [7:0] _seach_blockx_79_data_out;
  wire _seach_blockx_79_in_do;
  wire _seach_blockx_79_p_reset;
  wire _seach_blockx_79_m_clock;
  wire [7:0] _seach_blockx_78_map_block;
  wire [7:0] _seach_blockx_78_now;
  wire [7:0] _seach_blockx_78_start;
  wire [7:0] _seach_blockx_78_goal;
  wire [7:0] _seach_blockx_78_data_out;
  wire _seach_blockx_78_in_do;
  wire _seach_blockx_78_p_reset;
  wire _seach_blockx_78_m_clock;
  wire [7:0] _seach_blockx_77_map_block;
  wire [7:0] _seach_blockx_77_now;
  wire [7:0] _seach_blockx_77_start;
  wire [7:0] _seach_blockx_77_goal;
  wire [7:0] _seach_blockx_77_data_out;
  wire _seach_blockx_77_in_do;
  wire _seach_blockx_77_p_reset;
  wire _seach_blockx_77_m_clock;
  wire [7:0] _seach_blockx_76_map_block;
  wire [7:0] _seach_blockx_76_now;
  wire [7:0] _seach_blockx_76_start;
  wire [7:0] _seach_blockx_76_goal;
  wire [7:0] _seach_blockx_76_data_out;
  wire _seach_blockx_76_in_do;
  wire _seach_blockx_76_p_reset;
  wire _seach_blockx_76_m_clock;
  wire [7:0] _seach_blockx_75_map_block;
  wire [7:0] _seach_blockx_75_now;
  wire [7:0] _seach_blockx_75_start;
  wire [7:0] _seach_blockx_75_goal;
  wire [7:0] _seach_blockx_75_data_out;
  wire _seach_blockx_75_in_do;
  wire _seach_blockx_75_p_reset;
  wire _seach_blockx_75_m_clock;
  wire [7:0] _seach_blockx_74_map_block;
  wire [7:0] _seach_blockx_74_now;
  wire [7:0] _seach_blockx_74_start;
  wire [7:0] _seach_blockx_74_goal;
  wire [7:0] _seach_blockx_74_data_out;
  wire _seach_blockx_74_in_do;
  wire _seach_blockx_74_p_reset;
  wire _seach_blockx_74_m_clock;
  wire [7:0] _seach_blockx_73_map_block;
  wire [7:0] _seach_blockx_73_now;
  wire [7:0] _seach_blockx_73_start;
  wire [7:0] _seach_blockx_73_goal;
  wire [7:0] _seach_blockx_73_data_out;
  wire _seach_blockx_73_in_do;
  wire _seach_blockx_73_p_reset;
  wire _seach_blockx_73_m_clock;
  wire [7:0] _seach_blockx_72_map_block;
  wire [7:0] _seach_blockx_72_now;
  wire [7:0] _seach_blockx_72_start;
  wire [7:0] _seach_blockx_72_goal;
  wire [7:0] _seach_blockx_72_data_out;
  wire _seach_blockx_72_in_do;
  wire _seach_blockx_72_p_reset;
  wire _seach_blockx_72_m_clock;
  wire [7:0] _seach_blockx_71_map_block;
  wire [7:0] _seach_blockx_71_now;
  wire [7:0] _seach_blockx_71_start;
  wire [7:0] _seach_blockx_71_goal;
  wire [7:0] _seach_blockx_71_data_out;
  wire _seach_blockx_71_in_do;
  wire _seach_blockx_71_p_reset;
  wire _seach_blockx_71_m_clock;
  wire [7:0] _seach_blockx_70_map_block;
  wire [7:0] _seach_blockx_70_now;
  wire [7:0] _seach_blockx_70_start;
  wire [7:0] _seach_blockx_70_goal;
  wire [7:0] _seach_blockx_70_data_out;
  wire _seach_blockx_70_in_do;
  wire _seach_blockx_70_p_reset;
  wire _seach_blockx_70_m_clock;
  wire [7:0] _seach_blockx_69_map_block;
  wire [7:0] _seach_blockx_69_now;
  wire [7:0] _seach_blockx_69_start;
  wire [7:0] _seach_blockx_69_goal;
  wire [7:0] _seach_blockx_69_data_out;
  wire _seach_blockx_69_in_do;
  wire _seach_blockx_69_p_reset;
  wire _seach_blockx_69_m_clock;
  wire [7:0] _seach_blockx_68_map_block;
  wire [7:0] _seach_blockx_68_now;
  wire [7:0] _seach_blockx_68_start;
  wire [7:0] _seach_blockx_68_goal;
  wire [7:0] _seach_blockx_68_data_out;
  wire _seach_blockx_68_in_do;
  wire _seach_blockx_68_p_reset;
  wire _seach_blockx_68_m_clock;
  wire [7:0] _seach_blockx_67_map_block;
  wire [7:0] _seach_blockx_67_now;
  wire [7:0] _seach_blockx_67_start;
  wire [7:0] _seach_blockx_67_goal;
  wire [7:0] _seach_blockx_67_data_out;
  wire _seach_blockx_67_in_do;
  wire _seach_blockx_67_p_reset;
  wire _seach_blockx_67_m_clock;
  wire [7:0] _seach_blockx_66_map_block;
  wire [7:0] _seach_blockx_66_now;
  wire [7:0] _seach_blockx_66_start;
  wire [7:0] _seach_blockx_66_goal;
  wire [7:0] _seach_blockx_66_data_out;
  wire _seach_blockx_66_in_do;
  wire _seach_blockx_66_p_reset;
  wire _seach_blockx_66_m_clock;
  wire [7:0] _seach_blockx_65_map_block;
  wire [7:0] _seach_blockx_65_now;
  wire [7:0] _seach_blockx_65_start;
  wire [7:0] _seach_blockx_65_goal;
  wire [7:0] _seach_blockx_65_data_out;
  wire _seach_blockx_65_in_do;
  wire _seach_blockx_65_p_reset;
  wire _seach_blockx_65_m_clock;
  wire [7:0] _seach_blockx_64_map_block;
  wire [7:0] _seach_blockx_64_now;
  wire [7:0] _seach_blockx_64_start;
  wire [7:0] _seach_blockx_64_goal;
  wire [7:0] _seach_blockx_64_data_out;
  wire _seach_blockx_64_in_do;
  wire _seach_blockx_64_p_reset;
  wire _seach_blockx_64_m_clock;
  wire [7:0] _seach_blockx_63_map_block;
  wire [7:0] _seach_blockx_63_now;
  wire [7:0] _seach_blockx_63_start;
  wire [7:0] _seach_blockx_63_goal;
  wire [7:0] _seach_blockx_63_data_out;
  wire _seach_blockx_63_in_do;
  wire _seach_blockx_63_p_reset;
  wire _seach_blockx_63_m_clock;
  wire [7:0] _seach_blockx_62_map_block;
  wire [7:0] _seach_blockx_62_now;
  wire [7:0] _seach_blockx_62_start;
  wire [7:0] _seach_blockx_62_goal;
  wire [7:0] _seach_blockx_62_data_out;
  wire _seach_blockx_62_in_do;
  wire _seach_blockx_62_p_reset;
  wire _seach_blockx_62_m_clock;
  wire [7:0] _seach_blockx_61_map_block;
  wire [7:0] _seach_blockx_61_now;
  wire [7:0] _seach_blockx_61_start;
  wire [7:0] _seach_blockx_61_goal;
  wire [7:0] _seach_blockx_61_data_out;
  wire _seach_blockx_61_in_do;
  wire _seach_blockx_61_p_reset;
  wire _seach_blockx_61_m_clock;
  wire [7:0] _seach_blockx_60_map_block;
  wire [7:0] _seach_blockx_60_now;
  wire [7:0] _seach_blockx_60_start;
  wire [7:0] _seach_blockx_60_goal;
  wire [7:0] _seach_blockx_60_data_out;
  wire _seach_blockx_60_in_do;
  wire _seach_blockx_60_p_reset;
  wire _seach_blockx_60_m_clock;
  wire [7:0] _seach_blockx_59_map_block;
  wire [7:0] _seach_blockx_59_now;
  wire [7:0] _seach_blockx_59_start;
  wire [7:0] _seach_blockx_59_goal;
  wire [7:0] _seach_blockx_59_data_out;
  wire _seach_blockx_59_in_do;
  wire _seach_blockx_59_p_reset;
  wire _seach_blockx_59_m_clock;
  wire [7:0] _seach_blockx_58_map_block;
  wire [7:0] _seach_blockx_58_now;
  wire [7:0] _seach_blockx_58_start;
  wire [7:0] _seach_blockx_58_goal;
  wire [7:0] _seach_blockx_58_data_out;
  wire _seach_blockx_58_in_do;
  wire _seach_blockx_58_p_reset;
  wire _seach_blockx_58_m_clock;
  wire [7:0] _seach_blockx_57_map_block;
  wire [7:0] _seach_blockx_57_now;
  wire [7:0] _seach_blockx_57_start;
  wire [7:0] _seach_blockx_57_goal;
  wire [7:0] _seach_blockx_57_data_out;
  wire _seach_blockx_57_in_do;
  wire _seach_blockx_57_p_reset;
  wire _seach_blockx_57_m_clock;
  wire [7:0] _seach_blockx_56_map_block;
  wire [7:0] _seach_blockx_56_now;
  wire [7:0] _seach_blockx_56_start;
  wire [7:0] _seach_blockx_56_goal;
  wire [7:0] _seach_blockx_56_data_out;
  wire _seach_blockx_56_in_do;
  wire _seach_blockx_56_p_reset;
  wire _seach_blockx_56_m_clock;
  wire [7:0] _seach_blockx_55_map_block;
  wire [7:0] _seach_blockx_55_now;
  wire [7:0] _seach_blockx_55_start;
  wire [7:0] _seach_blockx_55_goal;
  wire [7:0] _seach_blockx_55_data_out;
  wire _seach_blockx_55_in_do;
  wire _seach_blockx_55_p_reset;
  wire _seach_blockx_55_m_clock;
  wire [7:0] _seach_blockx_54_map_block;
  wire [7:0] _seach_blockx_54_now;
  wire [7:0] _seach_blockx_54_start;
  wire [7:0] _seach_blockx_54_goal;
  wire [7:0] _seach_blockx_54_data_out;
  wire _seach_blockx_54_in_do;
  wire _seach_blockx_54_p_reset;
  wire _seach_blockx_54_m_clock;
  wire [7:0] _seach_blockx_53_map_block;
  wire [7:0] _seach_blockx_53_now;
  wire [7:0] _seach_blockx_53_start;
  wire [7:0] _seach_blockx_53_goal;
  wire [7:0] _seach_blockx_53_data_out;
  wire _seach_blockx_53_in_do;
  wire _seach_blockx_53_p_reset;
  wire _seach_blockx_53_m_clock;
  wire [7:0] _seach_blockx_52_map_block;
  wire [7:0] _seach_blockx_52_now;
  wire [7:0] _seach_blockx_52_start;
  wire [7:0] _seach_blockx_52_goal;
  wire [7:0] _seach_blockx_52_data_out;
  wire _seach_blockx_52_in_do;
  wire _seach_blockx_52_p_reset;
  wire _seach_blockx_52_m_clock;
  wire [7:0] _seach_blockx_51_map_block;
  wire [7:0] _seach_blockx_51_now;
  wire [7:0] _seach_blockx_51_start;
  wire [7:0] _seach_blockx_51_goal;
  wire [7:0] _seach_blockx_51_data_out;
  wire _seach_blockx_51_in_do;
  wire _seach_blockx_51_p_reset;
  wire _seach_blockx_51_m_clock;
  wire [7:0] _seach_blockx_50_map_block;
  wire [7:0] _seach_blockx_50_now;
  wire [7:0] _seach_blockx_50_start;
  wire [7:0] _seach_blockx_50_goal;
  wire [7:0] _seach_blockx_50_data_out;
  wire _seach_blockx_50_in_do;
  wire _seach_blockx_50_p_reset;
  wire _seach_blockx_50_m_clock;
  wire [7:0] _seach_blockx_49_map_block;
  wire [7:0] _seach_blockx_49_now;
  wire [7:0] _seach_blockx_49_start;
  wire [7:0] _seach_blockx_49_goal;
  wire [7:0] _seach_blockx_49_data_out;
  wire _seach_blockx_49_in_do;
  wire _seach_blockx_49_p_reset;
  wire _seach_blockx_49_m_clock;
  wire [7:0] _seach_blockx_48_map_block;
  wire [7:0] _seach_blockx_48_now;
  wire [7:0] _seach_blockx_48_start;
  wire [7:0] _seach_blockx_48_goal;
  wire [7:0] _seach_blockx_48_data_out;
  wire _seach_blockx_48_in_do;
  wire _seach_blockx_48_p_reset;
  wire _seach_blockx_48_m_clock;
  wire [7:0] _seach_blockx_47_map_block;
  wire [7:0] _seach_blockx_47_now;
  wire [7:0] _seach_blockx_47_start;
  wire [7:0] _seach_blockx_47_goal;
  wire [7:0] _seach_blockx_47_data_out;
  wire _seach_blockx_47_in_do;
  wire _seach_blockx_47_p_reset;
  wire _seach_blockx_47_m_clock;
  wire [7:0] _seach_blockx_46_map_block;
  wire [7:0] _seach_blockx_46_now;
  wire [7:0] _seach_blockx_46_start;
  wire [7:0] _seach_blockx_46_goal;
  wire [7:0] _seach_blockx_46_data_out;
  wire _seach_blockx_46_in_do;
  wire _seach_blockx_46_p_reset;
  wire _seach_blockx_46_m_clock;
  wire [7:0] _seach_blockx_45_map_block;
  wire [7:0] _seach_blockx_45_now;
  wire [7:0] _seach_blockx_45_start;
  wire [7:0] _seach_blockx_45_goal;
  wire [7:0] _seach_blockx_45_data_out;
  wire _seach_blockx_45_in_do;
  wire _seach_blockx_45_p_reset;
  wire _seach_blockx_45_m_clock;
  wire [7:0] _seach_blockx_44_map_block;
  wire [7:0] _seach_blockx_44_now;
  wire [7:0] _seach_blockx_44_start;
  wire [7:0] _seach_blockx_44_goal;
  wire [7:0] _seach_blockx_44_data_out;
  wire _seach_blockx_44_in_do;
  wire _seach_blockx_44_p_reset;
  wire _seach_blockx_44_m_clock;
  wire [7:0] _seach_blockx_43_map_block;
  wire [7:0] _seach_blockx_43_now;
  wire [7:0] _seach_blockx_43_start;
  wire [7:0] _seach_blockx_43_goal;
  wire [7:0] _seach_blockx_43_data_out;
  wire _seach_blockx_43_in_do;
  wire _seach_blockx_43_p_reset;
  wire _seach_blockx_43_m_clock;
  wire [7:0] _seach_blockx_42_map_block;
  wire [7:0] _seach_blockx_42_now;
  wire [7:0] _seach_blockx_42_start;
  wire [7:0] _seach_blockx_42_goal;
  wire [7:0] _seach_blockx_42_data_out;
  wire _seach_blockx_42_in_do;
  wire _seach_blockx_42_p_reset;
  wire _seach_blockx_42_m_clock;
  wire [7:0] _seach_blockx_41_map_block;
  wire [7:0] _seach_blockx_41_now;
  wire [7:0] _seach_blockx_41_start;
  wire [7:0] _seach_blockx_41_goal;
  wire [7:0] _seach_blockx_41_data_out;
  wire _seach_blockx_41_in_do;
  wire _seach_blockx_41_p_reset;
  wire _seach_blockx_41_m_clock;
  wire [7:0] _seach_blockx_40_map_block;
  wire [7:0] _seach_blockx_40_now;
  wire [7:0] _seach_blockx_40_start;
  wire [7:0] _seach_blockx_40_goal;
  wire [7:0] _seach_blockx_40_data_out;
  wire _seach_blockx_40_in_do;
  wire _seach_blockx_40_p_reset;
  wire _seach_blockx_40_m_clock;
  wire [7:0] _seach_blockx_39_map_block;
  wire [7:0] _seach_blockx_39_now;
  wire [7:0] _seach_blockx_39_start;
  wire [7:0] _seach_blockx_39_goal;
  wire [7:0] _seach_blockx_39_data_out;
  wire _seach_blockx_39_in_do;
  wire _seach_blockx_39_p_reset;
  wire _seach_blockx_39_m_clock;
  wire [7:0] _seach_blockx_38_map_block;
  wire [7:0] _seach_blockx_38_now;
  wire [7:0] _seach_blockx_38_start;
  wire [7:0] _seach_blockx_38_goal;
  wire [7:0] _seach_blockx_38_data_out;
  wire _seach_blockx_38_in_do;
  wire _seach_blockx_38_p_reset;
  wire _seach_blockx_38_m_clock;
  wire [7:0] _seach_blockx_37_map_block;
  wire [7:0] _seach_blockx_37_now;
  wire [7:0] _seach_blockx_37_start;
  wire [7:0] _seach_blockx_37_goal;
  wire [7:0] _seach_blockx_37_data_out;
  wire _seach_blockx_37_in_do;
  wire _seach_blockx_37_p_reset;
  wire _seach_blockx_37_m_clock;
  wire [7:0] _seach_blockx_36_map_block;
  wire [7:0] _seach_blockx_36_now;
  wire [7:0] _seach_blockx_36_start;
  wire [7:0] _seach_blockx_36_goal;
  wire [7:0] _seach_blockx_36_data_out;
  wire _seach_blockx_36_in_do;
  wire _seach_blockx_36_p_reset;
  wire _seach_blockx_36_m_clock;
  wire [7:0] _seach_blockx_35_map_block;
  wire [7:0] _seach_blockx_35_now;
  wire [7:0] _seach_blockx_35_start;
  wire [7:0] _seach_blockx_35_goal;
  wire [7:0] _seach_blockx_35_data_out;
  wire _seach_blockx_35_in_do;
  wire _seach_blockx_35_p_reset;
  wire _seach_blockx_35_m_clock;
  wire [7:0] _seach_blockx_34_map_block;
  wire [7:0] _seach_blockx_34_now;
  wire [7:0] _seach_blockx_34_start;
  wire [7:0] _seach_blockx_34_goal;
  wire [7:0] _seach_blockx_34_data_out;
  wire _seach_blockx_34_in_do;
  wire _seach_blockx_34_p_reset;
  wire _seach_blockx_34_m_clock;
  wire [7:0] _seach_blockx_33_map_block;
  wire [7:0] _seach_blockx_33_now;
  wire [7:0] _seach_blockx_33_start;
  wire [7:0] _seach_blockx_33_goal;
  wire [7:0] _seach_blockx_33_data_out;
  wire _seach_blockx_33_in_do;
  wire _seach_blockx_33_p_reset;
  wire _seach_blockx_33_m_clock;
  wire [7:0] _seach_blockx_32_map_block;
  wire [7:0] _seach_blockx_32_now;
  wire [7:0] _seach_blockx_32_start;
  wire [7:0] _seach_blockx_32_goal;
  wire [7:0] _seach_blockx_32_data_out;
  wire _seach_blockx_32_in_do;
  wire _seach_blockx_32_p_reset;
  wire _seach_blockx_32_m_clock;
  wire [7:0] _seach_blockx_31_map_block;
  wire [7:0] _seach_blockx_31_now;
  wire [7:0] _seach_blockx_31_start;
  wire [7:0] _seach_blockx_31_goal;
  wire [7:0] _seach_blockx_31_data_out;
  wire _seach_blockx_31_in_do;
  wire _seach_blockx_31_p_reset;
  wire _seach_blockx_31_m_clock;
  wire [7:0] _seach_blockx_30_map_block;
  wire [7:0] _seach_blockx_30_now;
  wire [7:0] _seach_blockx_30_start;
  wire [7:0] _seach_blockx_30_goal;
  wire [7:0] _seach_blockx_30_data_out;
  wire _seach_blockx_30_in_do;
  wire _seach_blockx_30_p_reset;
  wire _seach_blockx_30_m_clock;
  wire [7:0] _seach_blockx_29_map_block;
  wire [7:0] _seach_blockx_29_now;
  wire [7:0] _seach_blockx_29_start;
  wire [7:0] _seach_blockx_29_goal;
  wire [7:0] _seach_blockx_29_data_out;
  wire _seach_blockx_29_in_do;
  wire _seach_blockx_29_p_reset;
  wire _seach_blockx_29_m_clock;
  wire [7:0] _seach_blockx_28_map_block;
  wire [7:0] _seach_blockx_28_now;
  wire [7:0] _seach_blockx_28_start;
  wire [7:0] _seach_blockx_28_goal;
  wire [7:0] _seach_blockx_28_data_out;
  wire _seach_blockx_28_in_do;
  wire _seach_blockx_28_p_reset;
  wire _seach_blockx_28_m_clock;
  wire [7:0] _seach_blockx_27_map_block;
  wire [7:0] _seach_blockx_27_now;
  wire [7:0] _seach_blockx_27_start;
  wire [7:0] _seach_blockx_27_goal;
  wire [7:0] _seach_blockx_27_data_out;
  wire _seach_blockx_27_in_do;
  wire _seach_blockx_27_p_reset;
  wire _seach_blockx_27_m_clock;
  wire [7:0] _seach_blockx_26_map_block;
  wire [7:0] _seach_blockx_26_now;
  wire [7:0] _seach_blockx_26_start;
  wire [7:0] _seach_blockx_26_goal;
  wire [7:0] _seach_blockx_26_data_out;
  wire _seach_blockx_26_in_do;
  wire _seach_blockx_26_p_reset;
  wire _seach_blockx_26_m_clock;
  wire [7:0] _seach_blockx_25_map_block;
  wire [7:0] _seach_blockx_25_now;
  wire [7:0] _seach_blockx_25_start;
  wire [7:0] _seach_blockx_25_goal;
  wire [7:0] _seach_blockx_25_data_out;
  wire _seach_blockx_25_in_do;
  wire _seach_blockx_25_p_reset;
  wire _seach_blockx_25_m_clock;
  wire [7:0] _seach_blockx_24_map_block;
  wire [7:0] _seach_blockx_24_now;
  wire [7:0] _seach_blockx_24_start;
  wire [7:0] _seach_blockx_24_goal;
  wire [7:0] _seach_blockx_24_data_out;
  wire _seach_blockx_24_in_do;
  wire _seach_blockx_24_p_reset;
  wire _seach_blockx_24_m_clock;
  wire [7:0] _seach_blockx_23_map_block;
  wire [7:0] _seach_blockx_23_now;
  wire [7:0] _seach_blockx_23_start;
  wire [7:0] _seach_blockx_23_goal;
  wire [7:0] _seach_blockx_23_data_out;
  wire _seach_blockx_23_in_do;
  wire _seach_blockx_23_p_reset;
  wire _seach_blockx_23_m_clock;
  wire [7:0] _seach_blockx_22_map_block;
  wire [7:0] _seach_blockx_22_now;
  wire [7:0] _seach_blockx_22_start;
  wire [7:0] _seach_blockx_22_goal;
  wire [7:0] _seach_blockx_22_data_out;
  wire _seach_blockx_22_in_do;
  wire _seach_blockx_22_p_reset;
  wire _seach_blockx_22_m_clock;
  wire [7:0] _seach_blockx_21_map_block;
  wire [7:0] _seach_blockx_21_now;
  wire [7:0] _seach_blockx_21_start;
  wire [7:0] _seach_blockx_21_goal;
  wire [7:0] _seach_blockx_21_data_out;
  wire _seach_blockx_21_in_do;
  wire _seach_blockx_21_p_reset;
  wire _seach_blockx_21_m_clock;
  wire [7:0] _seach_blockx_20_map_block;
  wire [7:0] _seach_blockx_20_now;
  wire [7:0] _seach_blockx_20_start;
  wire [7:0] _seach_blockx_20_goal;
  wire [7:0] _seach_blockx_20_data_out;
  wire _seach_blockx_20_in_do;
  wire _seach_blockx_20_p_reset;
  wire _seach_blockx_20_m_clock;
  wire [7:0] _seach_blockx_19_map_block;
  wire [7:0] _seach_blockx_19_now;
  wire [7:0] _seach_blockx_19_start;
  wire [7:0] _seach_blockx_19_goal;
  wire [7:0] _seach_blockx_19_data_out;
  wire _seach_blockx_19_in_do;
  wire _seach_blockx_19_p_reset;
  wire _seach_blockx_19_m_clock;
  wire [7:0] _seach_blockx_18_map_block;
  wire [7:0] _seach_blockx_18_now;
  wire [7:0] _seach_blockx_18_start;
  wire [7:0] _seach_blockx_18_goal;
  wire [7:0] _seach_blockx_18_data_out;
  wire _seach_blockx_18_in_do;
  wire _seach_blockx_18_p_reset;
  wire _seach_blockx_18_m_clock;
  wire [7:0] _seach_blockx_17_map_block;
  wire [7:0] _seach_blockx_17_now;
  wire [7:0] _seach_blockx_17_start;
  wire [7:0] _seach_blockx_17_goal;
  wire [7:0] _seach_blockx_17_data_out;
  wire _seach_blockx_17_in_do;
  wire _seach_blockx_17_p_reset;
  wire _seach_blockx_17_m_clock;
  wire [7:0] _seach_blockx_16_map_block;
  wire [7:0] _seach_blockx_16_now;
  wire [7:0] _seach_blockx_16_start;
  wire [7:0] _seach_blockx_16_goal;
  wire [7:0] _seach_blockx_16_data_out;
  wire _seach_blockx_16_in_do;
  wire _seach_blockx_16_p_reset;
  wire _seach_blockx_16_m_clock;
  wire [7:0] _seach_blockx_15_map_block;
  wire [7:0] _seach_blockx_15_now;
  wire [7:0] _seach_blockx_15_start;
  wire [7:0] _seach_blockx_15_goal;
  wire [7:0] _seach_blockx_15_data_out;
  wire _seach_blockx_15_in_do;
  wire _seach_blockx_15_p_reset;
  wire _seach_blockx_15_m_clock;
  wire [7:0] _seach_blockx_14_map_block;
  wire [7:0] _seach_blockx_14_now;
  wire [7:0] _seach_blockx_14_start;
  wire [7:0] _seach_blockx_14_goal;
  wire [7:0] _seach_blockx_14_data_out;
  wire _seach_blockx_14_in_do;
  wire _seach_blockx_14_p_reset;
  wire _seach_blockx_14_m_clock;
  wire [7:0] _seach_blockx_13_map_block;
  wire [7:0] _seach_blockx_13_now;
  wire [7:0] _seach_blockx_13_start;
  wire [7:0] _seach_blockx_13_goal;
  wire [7:0] _seach_blockx_13_data_out;
  wire _seach_blockx_13_in_do;
  wire _seach_blockx_13_p_reset;
  wire _seach_blockx_13_m_clock;
  wire [7:0] _seach_blockx_12_map_block;
  wire [7:0] _seach_blockx_12_now;
  wire [7:0] _seach_blockx_12_start;
  wire [7:0] _seach_blockx_12_goal;
  wire [7:0] _seach_blockx_12_data_out;
  wire _seach_blockx_12_in_do;
  wire _seach_blockx_12_p_reset;
  wire _seach_blockx_12_m_clock;
  wire [7:0] _seach_blockx_11_map_block;
  wire [7:0] _seach_blockx_11_now;
  wire [7:0] _seach_blockx_11_start;
  wire [7:0] _seach_blockx_11_goal;
  wire [7:0] _seach_blockx_11_data_out;
  wire _seach_blockx_11_in_do;
  wire _seach_blockx_11_p_reset;
  wire _seach_blockx_11_m_clock;
  wire [7:0] _seach_blockx_10_map_block;
  wire [7:0] _seach_blockx_10_now;
  wire [7:0] _seach_blockx_10_start;
  wire [7:0] _seach_blockx_10_goal;
  wire [7:0] _seach_blockx_10_data_out;
  wire _seach_blockx_10_in_do;
  wire _seach_blockx_10_p_reset;
  wire _seach_blockx_10_m_clock;
  wire [7:0] _seach_blockx_9_map_block;
  wire [7:0] _seach_blockx_9_now;
  wire [7:0] _seach_blockx_9_start;
  wire [7:0] _seach_blockx_9_goal;
  wire [7:0] _seach_blockx_9_data_out;
  wire _seach_blockx_9_in_do;
  wire _seach_blockx_9_p_reset;
  wire _seach_blockx_9_m_clock;
  wire [7:0] _seach_blockx_8_map_block;
  wire [7:0] _seach_blockx_8_now;
  wire [7:0] _seach_blockx_8_start;
  wire [7:0] _seach_blockx_8_goal;
  wire [7:0] _seach_blockx_8_data_out;
  wire _seach_blockx_8_in_do;
  wire _seach_blockx_8_p_reset;
  wire _seach_blockx_8_m_clock;
  wire [7:0] _seach_blockx_7_map_block;
  wire [7:0] _seach_blockx_7_now;
  wire [7:0] _seach_blockx_7_start;
  wire [7:0] _seach_blockx_7_goal;
  wire [7:0] _seach_blockx_7_data_out;
  wire _seach_blockx_7_in_do;
  wire _seach_blockx_7_p_reset;
  wire _seach_blockx_7_m_clock;
  wire [7:0] _seach_blockx_6_map_block;
  wire [7:0] _seach_blockx_6_now;
  wire [7:0] _seach_blockx_6_start;
  wire [7:0] _seach_blockx_6_goal;
  wire [7:0] _seach_blockx_6_data_out;
  wire _seach_blockx_6_in_do;
  wire _seach_blockx_6_p_reset;
  wire _seach_blockx_6_m_clock;
  wire [7:0] _seach_blockx_5_map_block;
  wire [7:0] _seach_blockx_5_now;
  wire [7:0] _seach_blockx_5_start;
  wire [7:0] _seach_blockx_5_goal;
  wire [7:0] _seach_blockx_5_data_out;
  wire _seach_blockx_5_in_do;
  wire _seach_blockx_5_p_reset;
  wire _seach_blockx_5_m_clock;
  wire [7:0] _seach_blockx_4_map_block;
  wire [7:0] _seach_blockx_4_now;
  wire [7:0] _seach_blockx_4_start;
  wire [7:0] _seach_blockx_4_goal;
  wire [7:0] _seach_blockx_4_data_out;
  wire _seach_blockx_4_in_do;
  wire _seach_blockx_4_p_reset;
  wire _seach_blockx_4_m_clock;
  wire [7:0] _seach_blockx_3_map_block;
  wire [7:0] _seach_blockx_3_now;
  wire [7:0] _seach_blockx_3_start;
  wire [7:0] _seach_blockx_3_goal;
  wire [7:0] _seach_blockx_3_data_out;
  wire _seach_blockx_3_in_do;
  wire _seach_blockx_3_p_reset;
  wire _seach_blockx_3_m_clock;
  wire [7:0] _seach_blockx_2_map_block;
  wire [7:0] _seach_blockx_2_now;
  wire [7:0] _seach_blockx_2_start;
  wire [7:0] _seach_blockx_2_goal;
  wire [7:0] _seach_blockx_2_data_out;
  wire _seach_blockx_2_in_do;
  wire _seach_blockx_2_p_reset;
  wire _seach_blockx_2_m_clock;
  wire [7:0] _seach_blockx_1_map_block;
  wire [7:0] _seach_blockx_1_now;
  wire [7:0] _seach_blockx_1_start;
  wire [7:0] _seach_blockx_1_goal;
  wire [7:0] _seach_blockx_1_data_out;
  wire _seach_blockx_1_in_do;
  wire _seach_blockx_1_p_reset;
  wire _seach_blockx_1_m_clock;
  reg _reg_0;
  reg _reg_1;
seach_block seach_blockx (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_in_do), .start(_seach_blockx_start), .goal(_seach_blockx_goal), .data_out(_seach_blockx_data_out), .map_block(_seach_blockx_map_block), .now(_seach_blockx_now));
seach_block seach_blockx_195 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_195_in_do), .start(_seach_blockx_195_start), .goal(_seach_blockx_195_goal), .data_out(_seach_blockx_195_data_out), .map_block(_seach_blockx_195_map_block), .now(_seach_blockx_195_now));
seach_block seach_blockx_194 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_194_in_do), .start(_seach_blockx_194_start), .goal(_seach_blockx_194_goal), .data_out(_seach_blockx_194_data_out), .map_block(_seach_blockx_194_map_block), .now(_seach_blockx_194_now));
seach_block seach_blockx_193 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_193_in_do), .start(_seach_blockx_193_start), .goal(_seach_blockx_193_goal), .data_out(_seach_blockx_193_data_out), .map_block(_seach_blockx_193_map_block), .now(_seach_blockx_193_now));
seach_block seach_blockx_192 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_192_in_do), .start(_seach_blockx_192_start), .goal(_seach_blockx_192_goal), .data_out(_seach_blockx_192_data_out), .map_block(_seach_blockx_192_map_block), .now(_seach_blockx_192_now));
seach_block seach_blockx_191 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_191_in_do), .start(_seach_blockx_191_start), .goal(_seach_blockx_191_goal), .data_out(_seach_blockx_191_data_out), .map_block(_seach_blockx_191_map_block), .now(_seach_blockx_191_now));
seach_block seach_blockx_190 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_190_in_do), .start(_seach_blockx_190_start), .goal(_seach_blockx_190_goal), .data_out(_seach_blockx_190_data_out), .map_block(_seach_blockx_190_map_block), .now(_seach_blockx_190_now));
seach_block seach_blockx_189 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_189_in_do), .start(_seach_blockx_189_start), .goal(_seach_blockx_189_goal), .data_out(_seach_blockx_189_data_out), .map_block(_seach_blockx_189_map_block), .now(_seach_blockx_189_now));
seach_block seach_blockx_188 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_188_in_do), .start(_seach_blockx_188_start), .goal(_seach_blockx_188_goal), .data_out(_seach_blockx_188_data_out), .map_block(_seach_blockx_188_map_block), .now(_seach_blockx_188_now));
seach_block seach_blockx_187 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_187_in_do), .start(_seach_blockx_187_start), .goal(_seach_blockx_187_goal), .data_out(_seach_blockx_187_data_out), .map_block(_seach_blockx_187_map_block), .now(_seach_blockx_187_now));
seach_block seach_blockx_186 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_186_in_do), .start(_seach_blockx_186_start), .goal(_seach_blockx_186_goal), .data_out(_seach_blockx_186_data_out), .map_block(_seach_blockx_186_map_block), .now(_seach_blockx_186_now));
seach_block seach_blockx_185 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_185_in_do), .start(_seach_blockx_185_start), .goal(_seach_blockx_185_goal), .data_out(_seach_blockx_185_data_out), .map_block(_seach_blockx_185_map_block), .now(_seach_blockx_185_now));
seach_block seach_blockx_184 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_184_in_do), .start(_seach_blockx_184_start), .goal(_seach_blockx_184_goal), .data_out(_seach_blockx_184_data_out), .map_block(_seach_blockx_184_map_block), .now(_seach_blockx_184_now));
seach_block seach_blockx_183 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_183_in_do), .start(_seach_blockx_183_start), .goal(_seach_blockx_183_goal), .data_out(_seach_blockx_183_data_out), .map_block(_seach_blockx_183_map_block), .now(_seach_blockx_183_now));
seach_block seach_blockx_182 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_182_in_do), .start(_seach_blockx_182_start), .goal(_seach_blockx_182_goal), .data_out(_seach_blockx_182_data_out), .map_block(_seach_blockx_182_map_block), .now(_seach_blockx_182_now));
seach_block seach_blockx_181 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_181_in_do), .start(_seach_blockx_181_start), .goal(_seach_blockx_181_goal), .data_out(_seach_blockx_181_data_out), .map_block(_seach_blockx_181_map_block), .now(_seach_blockx_181_now));
seach_block seach_blockx_180 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_180_in_do), .start(_seach_blockx_180_start), .goal(_seach_blockx_180_goal), .data_out(_seach_blockx_180_data_out), .map_block(_seach_blockx_180_map_block), .now(_seach_blockx_180_now));
seach_block seach_blockx_179 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_179_in_do), .start(_seach_blockx_179_start), .goal(_seach_blockx_179_goal), .data_out(_seach_blockx_179_data_out), .map_block(_seach_blockx_179_map_block), .now(_seach_blockx_179_now));
seach_block seach_blockx_178 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_178_in_do), .start(_seach_blockx_178_start), .goal(_seach_blockx_178_goal), .data_out(_seach_blockx_178_data_out), .map_block(_seach_blockx_178_map_block), .now(_seach_blockx_178_now));
seach_block seach_blockx_177 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_177_in_do), .start(_seach_blockx_177_start), .goal(_seach_blockx_177_goal), .data_out(_seach_blockx_177_data_out), .map_block(_seach_blockx_177_map_block), .now(_seach_blockx_177_now));
seach_block seach_blockx_176 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_176_in_do), .start(_seach_blockx_176_start), .goal(_seach_blockx_176_goal), .data_out(_seach_blockx_176_data_out), .map_block(_seach_blockx_176_map_block), .now(_seach_blockx_176_now));
seach_block seach_blockx_175 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_175_in_do), .start(_seach_blockx_175_start), .goal(_seach_blockx_175_goal), .data_out(_seach_blockx_175_data_out), .map_block(_seach_blockx_175_map_block), .now(_seach_blockx_175_now));
seach_block seach_blockx_174 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_174_in_do), .start(_seach_blockx_174_start), .goal(_seach_blockx_174_goal), .data_out(_seach_blockx_174_data_out), .map_block(_seach_blockx_174_map_block), .now(_seach_blockx_174_now));
seach_block seach_blockx_173 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_173_in_do), .start(_seach_blockx_173_start), .goal(_seach_blockx_173_goal), .data_out(_seach_blockx_173_data_out), .map_block(_seach_blockx_173_map_block), .now(_seach_blockx_173_now));
seach_block seach_blockx_172 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_172_in_do), .start(_seach_blockx_172_start), .goal(_seach_blockx_172_goal), .data_out(_seach_blockx_172_data_out), .map_block(_seach_blockx_172_map_block), .now(_seach_blockx_172_now));
seach_block seach_blockx_171 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_171_in_do), .start(_seach_blockx_171_start), .goal(_seach_blockx_171_goal), .data_out(_seach_blockx_171_data_out), .map_block(_seach_blockx_171_map_block), .now(_seach_blockx_171_now));
seach_block seach_blockx_170 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_170_in_do), .start(_seach_blockx_170_start), .goal(_seach_blockx_170_goal), .data_out(_seach_blockx_170_data_out), .map_block(_seach_blockx_170_map_block), .now(_seach_blockx_170_now));
seach_block seach_blockx_169 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_169_in_do), .start(_seach_blockx_169_start), .goal(_seach_blockx_169_goal), .data_out(_seach_blockx_169_data_out), .map_block(_seach_blockx_169_map_block), .now(_seach_blockx_169_now));
seach_block seach_blockx_168 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_168_in_do), .start(_seach_blockx_168_start), .goal(_seach_blockx_168_goal), .data_out(_seach_blockx_168_data_out), .map_block(_seach_blockx_168_map_block), .now(_seach_blockx_168_now));
seach_block seach_blockx_167 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_167_in_do), .start(_seach_blockx_167_start), .goal(_seach_blockx_167_goal), .data_out(_seach_blockx_167_data_out), .map_block(_seach_blockx_167_map_block), .now(_seach_blockx_167_now));
seach_block seach_blockx_166 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_166_in_do), .start(_seach_blockx_166_start), .goal(_seach_blockx_166_goal), .data_out(_seach_blockx_166_data_out), .map_block(_seach_blockx_166_map_block), .now(_seach_blockx_166_now));
seach_block seach_blockx_165 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_165_in_do), .start(_seach_blockx_165_start), .goal(_seach_blockx_165_goal), .data_out(_seach_blockx_165_data_out), .map_block(_seach_blockx_165_map_block), .now(_seach_blockx_165_now));
seach_block seach_blockx_164 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_164_in_do), .start(_seach_blockx_164_start), .goal(_seach_blockx_164_goal), .data_out(_seach_blockx_164_data_out), .map_block(_seach_blockx_164_map_block), .now(_seach_blockx_164_now));
seach_block seach_blockx_163 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_163_in_do), .start(_seach_blockx_163_start), .goal(_seach_blockx_163_goal), .data_out(_seach_blockx_163_data_out), .map_block(_seach_blockx_163_map_block), .now(_seach_blockx_163_now));
seach_block seach_blockx_162 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_162_in_do), .start(_seach_blockx_162_start), .goal(_seach_blockx_162_goal), .data_out(_seach_blockx_162_data_out), .map_block(_seach_blockx_162_map_block), .now(_seach_blockx_162_now));
seach_block seach_blockx_161 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_161_in_do), .start(_seach_blockx_161_start), .goal(_seach_blockx_161_goal), .data_out(_seach_blockx_161_data_out), .map_block(_seach_blockx_161_map_block), .now(_seach_blockx_161_now));
seach_block seach_blockx_160 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_160_in_do), .start(_seach_blockx_160_start), .goal(_seach_blockx_160_goal), .data_out(_seach_blockx_160_data_out), .map_block(_seach_blockx_160_map_block), .now(_seach_blockx_160_now));
seach_block seach_blockx_159 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_159_in_do), .start(_seach_blockx_159_start), .goal(_seach_blockx_159_goal), .data_out(_seach_blockx_159_data_out), .map_block(_seach_blockx_159_map_block), .now(_seach_blockx_159_now));
seach_block seach_blockx_158 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_158_in_do), .start(_seach_blockx_158_start), .goal(_seach_blockx_158_goal), .data_out(_seach_blockx_158_data_out), .map_block(_seach_blockx_158_map_block), .now(_seach_blockx_158_now));
seach_block seach_blockx_157 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_157_in_do), .start(_seach_blockx_157_start), .goal(_seach_blockx_157_goal), .data_out(_seach_blockx_157_data_out), .map_block(_seach_blockx_157_map_block), .now(_seach_blockx_157_now));
seach_block seach_blockx_156 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_156_in_do), .start(_seach_blockx_156_start), .goal(_seach_blockx_156_goal), .data_out(_seach_blockx_156_data_out), .map_block(_seach_blockx_156_map_block), .now(_seach_blockx_156_now));
seach_block seach_blockx_155 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_155_in_do), .start(_seach_blockx_155_start), .goal(_seach_blockx_155_goal), .data_out(_seach_blockx_155_data_out), .map_block(_seach_blockx_155_map_block), .now(_seach_blockx_155_now));
seach_block seach_blockx_154 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_154_in_do), .start(_seach_blockx_154_start), .goal(_seach_blockx_154_goal), .data_out(_seach_blockx_154_data_out), .map_block(_seach_blockx_154_map_block), .now(_seach_blockx_154_now));
seach_block seach_blockx_153 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_153_in_do), .start(_seach_blockx_153_start), .goal(_seach_blockx_153_goal), .data_out(_seach_blockx_153_data_out), .map_block(_seach_blockx_153_map_block), .now(_seach_blockx_153_now));
seach_block seach_blockx_152 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_152_in_do), .start(_seach_blockx_152_start), .goal(_seach_blockx_152_goal), .data_out(_seach_blockx_152_data_out), .map_block(_seach_blockx_152_map_block), .now(_seach_blockx_152_now));
seach_block seach_blockx_151 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_151_in_do), .start(_seach_blockx_151_start), .goal(_seach_blockx_151_goal), .data_out(_seach_blockx_151_data_out), .map_block(_seach_blockx_151_map_block), .now(_seach_blockx_151_now));
seach_block seach_blockx_150 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_150_in_do), .start(_seach_blockx_150_start), .goal(_seach_blockx_150_goal), .data_out(_seach_blockx_150_data_out), .map_block(_seach_blockx_150_map_block), .now(_seach_blockx_150_now));
seach_block seach_blockx_149 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_149_in_do), .start(_seach_blockx_149_start), .goal(_seach_blockx_149_goal), .data_out(_seach_blockx_149_data_out), .map_block(_seach_blockx_149_map_block), .now(_seach_blockx_149_now));
seach_block seach_blockx_148 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_148_in_do), .start(_seach_blockx_148_start), .goal(_seach_blockx_148_goal), .data_out(_seach_blockx_148_data_out), .map_block(_seach_blockx_148_map_block), .now(_seach_blockx_148_now));
seach_block seach_blockx_147 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_147_in_do), .start(_seach_blockx_147_start), .goal(_seach_blockx_147_goal), .data_out(_seach_blockx_147_data_out), .map_block(_seach_blockx_147_map_block), .now(_seach_blockx_147_now));
seach_block seach_blockx_146 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_146_in_do), .start(_seach_blockx_146_start), .goal(_seach_blockx_146_goal), .data_out(_seach_blockx_146_data_out), .map_block(_seach_blockx_146_map_block), .now(_seach_blockx_146_now));
seach_block seach_blockx_145 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_145_in_do), .start(_seach_blockx_145_start), .goal(_seach_blockx_145_goal), .data_out(_seach_blockx_145_data_out), .map_block(_seach_blockx_145_map_block), .now(_seach_blockx_145_now));
seach_block seach_blockx_144 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_144_in_do), .start(_seach_blockx_144_start), .goal(_seach_blockx_144_goal), .data_out(_seach_blockx_144_data_out), .map_block(_seach_blockx_144_map_block), .now(_seach_blockx_144_now));
seach_block seach_blockx_143 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_143_in_do), .start(_seach_blockx_143_start), .goal(_seach_blockx_143_goal), .data_out(_seach_blockx_143_data_out), .map_block(_seach_blockx_143_map_block), .now(_seach_blockx_143_now));
seach_block seach_blockx_142 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_142_in_do), .start(_seach_blockx_142_start), .goal(_seach_blockx_142_goal), .data_out(_seach_blockx_142_data_out), .map_block(_seach_blockx_142_map_block), .now(_seach_blockx_142_now));
seach_block seach_blockx_141 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_141_in_do), .start(_seach_blockx_141_start), .goal(_seach_blockx_141_goal), .data_out(_seach_blockx_141_data_out), .map_block(_seach_blockx_141_map_block), .now(_seach_blockx_141_now));
seach_block seach_blockx_140 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_140_in_do), .start(_seach_blockx_140_start), .goal(_seach_blockx_140_goal), .data_out(_seach_blockx_140_data_out), .map_block(_seach_blockx_140_map_block), .now(_seach_blockx_140_now));
seach_block seach_blockx_139 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_139_in_do), .start(_seach_blockx_139_start), .goal(_seach_blockx_139_goal), .data_out(_seach_blockx_139_data_out), .map_block(_seach_blockx_139_map_block), .now(_seach_blockx_139_now));
seach_block seach_blockx_138 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_138_in_do), .start(_seach_blockx_138_start), .goal(_seach_blockx_138_goal), .data_out(_seach_blockx_138_data_out), .map_block(_seach_blockx_138_map_block), .now(_seach_blockx_138_now));
seach_block seach_blockx_137 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_137_in_do), .start(_seach_blockx_137_start), .goal(_seach_blockx_137_goal), .data_out(_seach_blockx_137_data_out), .map_block(_seach_blockx_137_map_block), .now(_seach_blockx_137_now));
seach_block seach_blockx_136 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_136_in_do), .start(_seach_blockx_136_start), .goal(_seach_blockx_136_goal), .data_out(_seach_blockx_136_data_out), .map_block(_seach_blockx_136_map_block), .now(_seach_blockx_136_now));
seach_block seach_blockx_135 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_135_in_do), .start(_seach_blockx_135_start), .goal(_seach_blockx_135_goal), .data_out(_seach_blockx_135_data_out), .map_block(_seach_blockx_135_map_block), .now(_seach_blockx_135_now));
seach_block seach_blockx_134 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_134_in_do), .start(_seach_blockx_134_start), .goal(_seach_blockx_134_goal), .data_out(_seach_blockx_134_data_out), .map_block(_seach_blockx_134_map_block), .now(_seach_blockx_134_now));
seach_block seach_blockx_133 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_133_in_do), .start(_seach_blockx_133_start), .goal(_seach_blockx_133_goal), .data_out(_seach_blockx_133_data_out), .map_block(_seach_blockx_133_map_block), .now(_seach_blockx_133_now));
seach_block seach_blockx_132 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_132_in_do), .start(_seach_blockx_132_start), .goal(_seach_blockx_132_goal), .data_out(_seach_blockx_132_data_out), .map_block(_seach_blockx_132_map_block), .now(_seach_blockx_132_now));
seach_block seach_blockx_131 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_131_in_do), .start(_seach_blockx_131_start), .goal(_seach_blockx_131_goal), .data_out(_seach_blockx_131_data_out), .map_block(_seach_blockx_131_map_block), .now(_seach_blockx_131_now));
seach_block seach_blockx_130 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_130_in_do), .start(_seach_blockx_130_start), .goal(_seach_blockx_130_goal), .data_out(_seach_blockx_130_data_out), .map_block(_seach_blockx_130_map_block), .now(_seach_blockx_130_now));
seach_block seach_blockx_129 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_129_in_do), .start(_seach_blockx_129_start), .goal(_seach_blockx_129_goal), .data_out(_seach_blockx_129_data_out), .map_block(_seach_blockx_129_map_block), .now(_seach_blockx_129_now));
seach_block seach_blockx_128 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_128_in_do), .start(_seach_blockx_128_start), .goal(_seach_blockx_128_goal), .data_out(_seach_blockx_128_data_out), .map_block(_seach_blockx_128_map_block), .now(_seach_blockx_128_now));
seach_block seach_blockx_127 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_127_in_do), .start(_seach_blockx_127_start), .goal(_seach_blockx_127_goal), .data_out(_seach_blockx_127_data_out), .map_block(_seach_blockx_127_map_block), .now(_seach_blockx_127_now));
seach_block seach_blockx_126 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_126_in_do), .start(_seach_blockx_126_start), .goal(_seach_blockx_126_goal), .data_out(_seach_blockx_126_data_out), .map_block(_seach_blockx_126_map_block), .now(_seach_blockx_126_now));
seach_block seach_blockx_125 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_125_in_do), .start(_seach_blockx_125_start), .goal(_seach_blockx_125_goal), .data_out(_seach_blockx_125_data_out), .map_block(_seach_blockx_125_map_block), .now(_seach_blockx_125_now));
seach_block seach_blockx_124 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_124_in_do), .start(_seach_blockx_124_start), .goal(_seach_blockx_124_goal), .data_out(_seach_blockx_124_data_out), .map_block(_seach_blockx_124_map_block), .now(_seach_blockx_124_now));
seach_block seach_blockx_123 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_123_in_do), .start(_seach_blockx_123_start), .goal(_seach_blockx_123_goal), .data_out(_seach_blockx_123_data_out), .map_block(_seach_blockx_123_map_block), .now(_seach_blockx_123_now));
seach_block seach_blockx_122 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_122_in_do), .start(_seach_blockx_122_start), .goal(_seach_blockx_122_goal), .data_out(_seach_blockx_122_data_out), .map_block(_seach_blockx_122_map_block), .now(_seach_blockx_122_now));
seach_block seach_blockx_121 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_121_in_do), .start(_seach_blockx_121_start), .goal(_seach_blockx_121_goal), .data_out(_seach_blockx_121_data_out), .map_block(_seach_blockx_121_map_block), .now(_seach_blockx_121_now));
seach_block seach_blockx_120 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_120_in_do), .start(_seach_blockx_120_start), .goal(_seach_blockx_120_goal), .data_out(_seach_blockx_120_data_out), .map_block(_seach_blockx_120_map_block), .now(_seach_blockx_120_now));
seach_block seach_blockx_119 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_119_in_do), .start(_seach_blockx_119_start), .goal(_seach_blockx_119_goal), .data_out(_seach_blockx_119_data_out), .map_block(_seach_blockx_119_map_block), .now(_seach_blockx_119_now));
seach_block seach_blockx_118 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_118_in_do), .start(_seach_blockx_118_start), .goal(_seach_blockx_118_goal), .data_out(_seach_blockx_118_data_out), .map_block(_seach_blockx_118_map_block), .now(_seach_blockx_118_now));
seach_block seach_blockx_117 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_117_in_do), .start(_seach_blockx_117_start), .goal(_seach_blockx_117_goal), .data_out(_seach_blockx_117_data_out), .map_block(_seach_blockx_117_map_block), .now(_seach_blockx_117_now));
seach_block seach_blockx_116 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_116_in_do), .start(_seach_blockx_116_start), .goal(_seach_blockx_116_goal), .data_out(_seach_blockx_116_data_out), .map_block(_seach_blockx_116_map_block), .now(_seach_blockx_116_now));
seach_block seach_blockx_115 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_115_in_do), .start(_seach_blockx_115_start), .goal(_seach_blockx_115_goal), .data_out(_seach_blockx_115_data_out), .map_block(_seach_blockx_115_map_block), .now(_seach_blockx_115_now));
seach_block seach_blockx_114 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_114_in_do), .start(_seach_blockx_114_start), .goal(_seach_blockx_114_goal), .data_out(_seach_blockx_114_data_out), .map_block(_seach_blockx_114_map_block), .now(_seach_blockx_114_now));
seach_block seach_blockx_113 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_113_in_do), .start(_seach_blockx_113_start), .goal(_seach_blockx_113_goal), .data_out(_seach_blockx_113_data_out), .map_block(_seach_blockx_113_map_block), .now(_seach_blockx_113_now));
seach_block seach_blockx_112 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_112_in_do), .start(_seach_blockx_112_start), .goal(_seach_blockx_112_goal), .data_out(_seach_blockx_112_data_out), .map_block(_seach_blockx_112_map_block), .now(_seach_blockx_112_now));
seach_block seach_blockx_111 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_111_in_do), .start(_seach_blockx_111_start), .goal(_seach_blockx_111_goal), .data_out(_seach_blockx_111_data_out), .map_block(_seach_blockx_111_map_block), .now(_seach_blockx_111_now));
seach_block seach_blockx_110 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_110_in_do), .start(_seach_blockx_110_start), .goal(_seach_blockx_110_goal), .data_out(_seach_blockx_110_data_out), .map_block(_seach_blockx_110_map_block), .now(_seach_blockx_110_now));
seach_block seach_blockx_109 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_109_in_do), .start(_seach_blockx_109_start), .goal(_seach_blockx_109_goal), .data_out(_seach_blockx_109_data_out), .map_block(_seach_blockx_109_map_block), .now(_seach_blockx_109_now));
seach_block seach_blockx_108 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_108_in_do), .start(_seach_blockx_108_start), .goal(_seach_blockx_108_goal), .data_out(_seach_blockx_108_data_out), .map_block(_seach_blockx_108_map_block), .now(_seach_blockx_108_now));
seach_block seach_blockx_107 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_107_in_do), .start(_seach_blockx_107_start), .goal(_seach_blockx_107_goal), .data_out(_seach_blockx_107_data_out), .map_block(_seach_blockx_107_map_block), .now(_seach_blockx_107_now));
seach_block seach_blockx_106 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_106_in_do), .start(_seach_blockx_106_start), .goal(_seach_blockx_106_goal), .data_out(_seach_blockx_106_data_out), .map_block(_seach_blockx_106_map_block), .now(_seach_blockx_106_now));
seach_block seach_blockx_105 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_105_in_do), .start(_seach_blockx_105_start), .goal(_seach_blockx_105_goal), .data_out(_seach_blockx_105_data_out), .map_block(_seach_blockx_105_map_block), .now(_seach_blockx_105_now));
seach_block seach_blockx_104 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_104_in_do), .start(_seach_blockx_104_start), .goal(_seach_blockx_104_goal), .data_out(_seach_blockx_104_data_out), .map_block(_seach_blockx_104_map_block), .now(_seach_blockx_104_now));
seach_block seach_blockx_103 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_103_in_do), .start(_seach_blockx_103_start), .goal(_seach_blockx_103_goal), .data_out(_seach_blockx_103_data_out), .map_block(_seach_blockx_103_map_block), .now(_seach_blockx_103_now));
seach_block seach_blockx_102 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_102_in_do), .start(_seach_blockx_102_start), .goal(_seach_blockx_102_goal), .data_out(_seach_blockx_102_data_out), .map_block(_seach_blockx_102_map_block), .now(_seach_blockx_102_now));
seach_block seach_blockx_101 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_101_in_do), .start(_seach_blockx_101_start), .goal(_seach_blockx_101_goal), .data_out(_seach_blockx_101_data_out), .map_block(_seach_blockx_101_map_block), .now(_seach_blockx_101_now));
seach_block seach_blockx_100 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_100_in_do), .start(_seach_blockx_100_start), .goal(_seach_blockx_100_goal), .data_out(_seach_blockx_100_data_out), .map_block(_seach_blockx_100_map_block), .now(_seach_blockx_100_now));
seach_block seach_blockx_99 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_99_in_do), .start(_seach_blockx_99_start), .goal(_seach_blockx_99_goal), .data_out(_seach_blockx_99_data_out), .map_block(_seach_blockx_99_map_block), .now(_seach_blockx_99_now));
seach_block seach_blockx_98 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_98_in_do), .start(_seach_blockx_98_start), .goal(_seach_blockx_98_goal), .data_out(_seach_blockx_98_data_out), .map_block(_seach_blockx_98_map_block), .now(_seach_blockx_98_now));
seach_block seach_blockx_97 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_97_in_do), .start(_seach_blockx_97_start), .goal(_seach_blockx_97_goal), .data_out(_seach_blockx_97_data_out), .map_block(_seach_blockx_97_map_block), .now(_seach_blockx_97_now));
seach_block seach_blockx_96 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_96_in_do), .start(_seach_blockx_96_start), .goal(_seach_blockx_96_goal), .data_out(_seach_blockx_96_data_out), .map_block(_seach_blockx_96_map_block), .now(_seach_blockx_96_now));
seach_block seach_blockx_95 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_95_in_do), .start(_seach_blockx_95_start), .goal(_seach_blockx_95_goal), .data_out(_seach_blockx_95_data_out), .map_block(_seach_blockx_95_map_block), .now(_seach_blockx_95_now));
seach_block seach_blockx_94 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_94_in_do), .start(_seach_blockx_94_start), .goal(_seach_blockx_94_goal), .data_out(_seach_blockx_94_data_out), .map_block(_seach_blockx_94_map_block), .now(_seach_blockx_94_now));
seach_block seach_blockx_93 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_93_in_do), .start(_seach_blockx_93_start), .goal(_seach_blockx_93_goal), .data_out(_seach_blockx_93_data_out), .map_block(_seach_blockx_93_map_block), .now(_seach_blockx_93_now));
seach_block seach_blockx_92 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_92_in_do), .start(_seach_blockx_92_start), .goal(_seach_blockx_92_goal), .data_out(_seach_blockx_92_data_out), .map_block(_seach_blockx_92_map_block), .now(_seach_blockx_92_now));
seach_block seach_blockx_91 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_91_in_do), .start(_seach_blockx_91_start), .goal(_seach_blockx_91_goal), .data_out(_seach_blockx_91_data_out), .map_block(_seach_blockx_91_map_block), .now(_seach_blockx_91_now));
seach_block seach_blockx_90 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_90_in_do), .start(_seach_blockx_90_start), .goal(_seach_blockx_90_goal), .data_out(_seach_blockx_90_data_out), .map_block(_seach_blockx_90_map_block), .now(_seach_blockx_90_now));
seach_block seach_blockx_89 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_89_in_do), .start(_seach_blockx_89_start), .goal(_seach_blockx_89_goal), .data_out(_seach_blockx_89_data_out), .map_block(_seach_blockx_89_map_block), .now(_seach_blockx_89_now));
seach_block seach_blockx_88 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_88_in_do), .start(_seach_blockx_88_start), .goal(_seach_blockx_88_goal), .data_out(_seach_blockx_88_data_out), .map_block(_seach_blockx_88_map_block), .now(_seach_blockx_88_now));
seach_block seach_blockx_87 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_87_in_do), .start(_seach_blockx_87_start), .goal(_seach_blockx_87_goal), .data_out(_seach_blockx_87_data_out), .map_block(_seach_blockx_87_map_block), .now(_seach_blockx_87_now));
seach_block seach_blockx_86 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_86_in_do), .start(_seach_blockx_86_start), .goal(_seach_blockx_86_goal), .data_out(_seach_blockx_86_data_out), .map_block(_seach_blockx_86_map_block), .now(_seach_blockx_86_now));
seach_block seach_blockx_85 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_85_in_do), .start(_seach_blockx_85_start), .goal(_seach_blockx_85_goal), .data_out(_seach_blockx_85_data_out), .map_block(_seach_blockx_85_map_block), .now(_seach_blockx_85_now));
seach_block seach_blockx_84 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_84_in_do), .start(_seach_blockx_84_start), .goal(_seach_blockx_84_goal), .data_out(_seach_blockx_84_data_out), .map_block(_seach_blockx_84_map_block), .now(_seach_blockx_84_now));
seach_block seach_blockx_83 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_83_in_do), .start(_seach_blockx_83_start), .goal(_seach_blockx_83_goal), .data_out(_seach_blockx_83_data_out), .map_block(_seach_blockx_83_map_block), .now(_seach_blockx_83_now));
seach_block seach_blockx_82 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_82_in_do), .start(_seach_blockx_82_start), .goal(_seach_blockx_82_goal), .data_out(_seach_blockx_82_data_out), .map_block(_seach_blockx_82_map_block), .now(_seach_blockx_82_now));
seach_block seach_blockx_81 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_81_in_do), .start(_seach_blockx_81_start), .goal(_seach_blockx_81_goal), .data_out(_seach_blockx_81_data_out), .map_block(_seach_blockx_81_map_block), .now(_seach_blockx_81_now));
seach_block seach_blockx_80 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_80_in_do), .start(_seach_blockx_80_start), .goal(_seach_blockx_80_goal), .data_out(_seach_blockx_80_data_out), .map_block(_seach_blockx_80_map_block), .now(_seach_blockx_80_now));
seach_block seach_blockx_79 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_79_in_do), .start(_seach_blockx_79_start), .goal(_seach_blockx_79_goal), .data_out(_seach_blockx_79_data_out), .map_block(_seach_blockx_79_map_block), .now(_seach_blockx_79_now));
seach_block seach_blockx_78 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_78_in_do), .start(_seach_blockx_78_start), .goal(_seach_blockx_78_goal), .data_out(_seach_blockx_78_data_out), .map_block(_seach_blockx_78_map_block), .now(_seach_blockx_78_now));
seach_block seach_blockx_77 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_77_in_do), .start(_seach_blockx_77_start), .goal(_seach_blockx_77_goal), .data_out(_seach_blockx_77_data_out), .map_block(_seach_blockx_77_map_block), .now(_seach_blockx_77_now));
seach_block seach_blockx_76 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_76_in_do), .start(_seach_blockx_76_start), .goal(_seach_blockx_76_goal), .data_out(_seach_blockx_76_data_out), .map_block(_seach_blockx_76_map_block), .now(_seach_blockx_76_now));
seach_block seach_blockx_75 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_75_in_do), .start(_seach_blockx_75_start), .goal(_seach_blockx_75_goal), .data_out(_seach_blockx_75_data_out), .map_block(_seach_blockx_75_map_block), .now(_seach_blockx_75_now));
seach_block seach_blockx_74 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_74_in_do), .start(_seach_blockx_74_start), .goal(_seach_blockx_74_goal), .data_out(_seach_blockx_74_data_out), .map_block(_seach_blockx_74_map_block), .now(_seach_blockx_74_now));
seach_block seach_blockx_73 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_73_in_do), .start(_seach_blockx_73_start), .goal(_seach_blockx_73_goal), .data_out(_seach_blockx_73_data_out), .map_block(_seach_blockx_73_map_block), .now(_seach_blockx_73_now));
seach_block seach_blockx_72 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_72_in_do), .start(_seach_blockx_72_start), .goal(_seach_blockx_72_goal), .data_out(_seach_blockx_72_data_out), .map_block(_seach_blockx_72_map_block), .now(_seach_blockx_72_now));
seach_block seach_blockx_71 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_71_in_do), .start(_seach_blockx_71_start), .goal(_seach_blockx_71_goal), .data_out(_seach_blockx_71_data_out), .map_block(_seach_blockx_71_map_block), .now(_seach_blockx_71_now));
seach_block seach_blockx_70 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_70_in_do), .start(_seach_blockx_70_start), .goal(_seach_blockx_70_goal), .data_out(_seach_blockx_70_data_out), .map_block(_seach_blockx_70_map_block), .now(_seach_blockx_70_now));
seach_block seach_blockx_69 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_69_in_do), .start(_seach_blockx_69_start), .goal(_seach_blockx_69_goal), .data_out(_seach_blockx_69_data_out), .map_block(_seach_blockx_69_map_block), .now(_seach_blockx_69_now));
seach_block seach_blockx_68 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_68_in_do), .start(_seach_blockx_68_start), .goal(_seach_blockx_68_goal), .data_out(_seach_blockx_68_data_out), .map_block(_seach_blockx_68_map_block), .now(_seach_blockx_68_now));
seach_block seach_blockx_67 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_67_in_do), .start(_seach_blockx_67_start), .goal(_seach_blockx_67_goal), .data_out(_seach_blockx_67_data_out), .map_block(_seach_blockx_67_map_block), .now(_seach_blockx_67_now));
seach_block seach_blockx_66 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_66_in_do), .start(_seach_blockx_66_start), .goal(_seach_blockx_66_goal), .data_out(_seach_blockx_66_data_out), .map_block(_seach_blockx_66_map_block), .now(_seach_blockx_66_now));
seach_block seach_blockx_65 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_65_in_do), .start(_seach_blockx_65_start), .goal(_seach_blockx_65_goal), .data_out(_seach_blockx_65_data_out), .map_block(_seach_blockx_65_map_block), .now(_seach_blockx_65_now));
seach_block seach_blockx_64 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_64_in_do), .start(_seach_blockx_64_start), .goal(_seach_blockx_64_goal), .data_out(_seach_blockx_64_data_out), .map_block(_seach_blockx_64_map_block), .now(_seach_blockx_64_now));
seach_block seach_blockx_63 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_63_in_do), .start(_seach_blockx_63_start), .goal(_seach_blockx_63_goal), .data_out(_seach_blockx_63_data_out), .map_block(_seach_blockx_63_map_block), .now(_seach_blockx_63_now));
seach_block seach_blockx_62 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_62_in_do), .start(_seach_blockx_62_start), .goal(_seach_blockx_62_goal), .data_out(_seach_blockx_62_data_out), .map_block(_seach_blockx_62_map_block), .now(_seach_blockx_62_now));
seach_block seach_blockx_61 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_61_in_do), .start(_seach_blockx_61_start), .goal(_seach_blockx_61_goal), .data_out(_seach_blockx_61_data_out), .map_block(_seach_blockx_61_map_block), .now(_seach_blockx_61_now));
seach_block seach_blockx_60 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_60_in_do), .start(_seach_blockx_60_start), .goal(_seach_blockx_60_goal), .data_out(_seach_blockx_60_data_out), .map_block(_seach_blockx_60_map_block), .now(_seach_blockx_60_now));
seach_block seach_blockx_59 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_59_in_do), .start(_seach_blockx_59_start), .goal(_seach_blockx_59_goal), .data_out(_seach_blockx_59_data_out), .map_block(_seach_blockx_59_map_block), .now(_seach_blockx_59_now));
seach_block seach_blockx_58 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_58_in_do), .start(_seach_blockx_58_start), .goal(_seach_blockx_58_goal), .data_out(_seach_blockx_58_data_out), .map_block(_seach_blockx_58_map_block), .now(_seach_blockx_58_now));
seach_block seach_blockx_57 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_57_in_do), .start(_seach_blockx_57_start), .goal(_seach_blockx_57_goal), .data_out(_seach_blockx_57_data_out), .map_block(_seach_blockx_57_map_block), .now(_seach_blockx_57_now));
seach_block seach_blockx_56 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_56_in_do), .start(_seach_blockx_56_start), .goal(_seach_blockx_56_goal), .data_out(_seach_blockx_56_data_out), .map_block(_seach_blockx_56_map_block), .now(_seach_blockx_56_now));
seach_block seach_blockx_55 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_55_in_do), .start(_seach_blockx_55_start), .goal(_seach_blockx_55_goal), .data_out(_seach_blockx_55_data_out), .map_block(_seach_blockx_55_map_block), .now(_seach_blockx_55_now));
seach_block seach_blockx_54 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_54_in_do), .start(_seach_blockx_54_start), .goal(_seach_blockx_54_goal), .data_out(_seach_blockx_54_data_out), .map_block(_seach_blockx_54_map_block), .now(_seach_blockx_54_now));
seach_block seach_blockx_53 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_53_in_do), .start(_seach_blockx_53_start), .goal(_seach_blockx_53_goal), .data_out(_seach_blockx_53_data_out), .map_block(_seach_blockx_53_map_block), .now(_seach_blockx_53_now));
seach_block seach_blockx_52 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_52_in_do), .start(_seach_blockx_52_start), .goal(_seach_blockx_52_goal), .data_out(_seach_blockx_52_data_out), .map_block(_seach_blockx_52_map_block), .now(_seach_blockx_52_now));
seach_block seach_blockx_51 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_51_in_do), .start(_seach_blockx_51_start), .goal(_seach_blockx_51_goal), .data_out(_seach_blockx_51_data_out), .map_block(_seach_blockx_51_map_block), .now(_seach_blockx_51_now));
seach_block seach_blockx_50 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_50_in_do), .start(_seach_blockx_50_start), .goal(_seach_blockx_50_goal), .data_out(_seach_blockx_50_data_out), .map_block(_seach_blockx_50_map_block), .now(_seach_blockx_50_now));
seach_block seach_blockx_49 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_49_in_do), .start(_seach_blockx_49_start), .goal(_seach_blockx_49_goal), .data_out(_seach_blockx_49_data_out), .map_block(_seach_blockx_49_map_block), .now(_seach_blockx_49_now));
seach_block seach_blockx_48 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_48_in_do), .start(_seach_blockx_48_start), .goal(_seach_blockx_48_goal), .data_out(_seach_blockx_48_data_out), .map_block(_seach_blockx_48_map_block), .now(_seach_blockx_48_now));
seach_block seach_blockx_47 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_47_in_do), .start(_seach_blockx_47_start), .goal(_seach_blockx_47_goal), .data_out(_seach_blockx_47_data_out), .map_block(_seach_blockx_47_map_block), .now(_seach_blockx_47_now));
seach_block seach_blockx_46 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_46_in_do), .start(_seach_blockx_46_start), .goal(_seach_blockx_46_goal), .data_out(_seach_blockx_46_data_out), .map_block(_seach_blockx_46_map_block), .now(_seach_blockx_46_now));
seach_block seach_blockx_45 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_45_in_do), .start(_seach_blockx_45_start), .goal(_seach_blockx_45_goal), .data_out(_seach_blockx_45_data_out), .map_block(_seach_blockx_45_map_block), .now(_seach_blockx_45_now));
seach_block seach_blockx_44 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_44_in_do), .start(_seach_blockx_44_start), .goal(_seach_blockx_44_goal), .data_out(_seach_blockx_44_data_out), .map_block(_seach_blockx_44_map_block), .now(_seach_blockx_44_now));
seach_block seach_blockx_43 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_43_in_do), .start(_seach_blockx_43_start), .goal(_seach_blockx_43_goal), .data_out(_seach_blockx_43_data_out), .map_block(_seach_blockx_43_map_block), .now(_seach_blockx_43_now));
seach_block seach_blockx_42 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_42_in_do), .start(_seach_blockx_42_start), .goal(_seach_blockx_42_goal), .data_out(_seach_blockx_42_data_out), .map_block(_seach_blockx_42_map_block), .now(_seach_blockx_42_now));
seach_block seach_blockx_41 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_41_in_do), .start(_seach_blockx_41_start), .goal(_seach_blockx_41_goal), .data_out(_seach_blockx_41_data_out), .map_block(_seach_blockx_41_map_block), .now(_seach_blockx_41_now));
seach_block seach_blockx_40 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_40_in_do), .start(_seach_blockx_40_start), .goal(_seach_blockx_40_goal), .data_out(_seach_blockx_40_data_out), .map_block(_seach_blockx_40_map_block), .now(_seach_blockx_40_now));
seach_block seach_blockx_39 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_39_in_do), .start(_seach_blockx_39_start), .goal(_seach_blockx_39_goal), .data_out(_seach_blockx_39_data_out), .map_block(_seach_blockx_39_map_block), .now(_seach_blockx_39_now));
seach_block seach_blockx_38 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_38_in_do), .start(_seach_blockx_38_start), .goal(_seach_blockx_38_goal), .data_out(_seach_blockx_38_data_out), .map_block(_seach_blockx_38_map_block), .now(_seach_blockx_38_now));
seach_block seach_blockx_37 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_37_in_do), .start(_seach_blockx_37_start), .goal(_seach_blockx_37_goal), .data_out(_seach_blockx_37_data_out), .map_block(_seach_blockx_37_map_block), .now(_seach_blockx_37_now));
seach_block seach_blockx_36 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_36_in_do), .start(_seach_blockx_36_start), .goal(_seach_blockx_36_goal), .data_out(_seach_blockx_36_data_out), .map_block(_seach_blockx_36_map_block), .now(_seach_blockx_36_now));
seach_block seach_blockx_35 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_35_in_do), .start(_seach_blockx_35_start), .goal(_seach_blockx_35_goal), .data_out(_seach_blockx_35_data_out), .map_block(_seach_blockx_35_map_block), .now(_seach_blockx_35_now));
seach_block seach_blockx_34 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_34_in_do), .start(_seach_blockx_34_start), .goal(_seach_blockx_34_goal), .data_out(_seach_blockx_34_data_out), .map_block(_seach_blockx_34_map_block), .now(_seach_blockx_34_now));
seach_block seach_blockx_33 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_33_in_do), .start(_seach_blockx_33_start), .goal(_seach_blockx_33_goal), .data_out(_seach_blockx_33_data_out), .map_block(_seach_blockx_33_map_block), .now(_seach_blockx_33_now));
seach_block seach_blockx_32 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_32_in_do), .start(_seach_blockx_32_start), .goal(_seach_blockx_32_goal), .data_out(_seach_blockx_32_data_out), .map_block(_seach_blockx_32_map_block), .now(_seach_blockx_32_now));
seach_block seach_blockx_31 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_31_in_do), .start(_seach_blockx_31_start), .goal(_seach_blockx_31_goal), .data_out(_seach_blockx_31_data_out), .map_block(_seach_blockx_31_map_block), .now(_seach_blockx_31_now));
seach_block seach_blockx_30 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_30_in_do), .start(_seach_blockx_30_start), .goal(_seach_blockx_30_goal), .data_out(_seach_blockx_30_data_out), .map_block(_seach_blockx_30_map_block), .now(_seach_blockx_30_now));
seach_block seach_blockx_29 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_29_in_do), .start(_seach_blockx_29_start), .goal(_seach_blockx_29_goal), .data_out(_seach_blockx_29_data_out), .map_block(_seach_blockx_29_map_block), .now(_seach_blockx_29_now));
seach_block seach_blockx_28 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_28_in_do), .start(_seach_blockx_28_start), .goal(_seach_blockx_28_goal), .data_out(_seach_blockx_28_data_out), .map_block(_seach_blockx_28_map_block), .now(_seach_blockx_28_now));
seach_block seach_blockx_27 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_27_in_do), .start(_seach_blockx_27_start), .goal(_seach_blockx_27_goal), .data_out(_seach_blockx_27_data_out), .map_block(_seach_blockx_27_map_block), .now(_seach_blockx_27_now));
seach_block seach_blockx_26 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_26_in_do), .start(_seach_blockx_26_start), .goal(_seach_blockx_26_goal), .data_out(_seach_blockx_26_data_out), .map_block(_seach_blockx_26_map_block), .now(_seach_blockx_26_now));
seach_block seach_blockx_25 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_25_in_do), .start(_seach_blockx_25_start), .goal(_seach_blockx_25_goal), .data_out(_seach_blockx_25_data_out), .map_block(_seach_blockx_25_map_block), .now(_seach_blockx_25_now));
seach_block seach_blockx_24 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_24_in_do), .start(_seach_blockx_24_start), .goal(_seach_blockx_24_goal), .data_out(_seach_blockx_24_data_out), .map_block(_seach_blockx_24_map_block), .now(_seach_blockx_24_now));
seach_block seach_blockx_23 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_23_in_do), .start(_seach_blockx_23_start), .goal(_seach_blockx_23_goal), .data_out(_seach_blockx_23_data_out), .map_block(_seach_blockx_23_map_block), .now(_seach_blockx_23_now));
seach_block seach_blockx_22 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_22_in_do), .start(_seach_blockx_22_start), .goal(_seach_blockx_22_goal), .data_out(_seach_blockx_22_data_out), .map_block(_seach_blockx_22_map_block), .now(_seach_blockx_22_now));
seach_block seach_blockx_21 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_21_in_do), .start(_seach_blockx_21_start), .goal(_seach_blockx_21_goal), .data_out(_seach_blockx_21_data_out), .map_block(_seach_blockx_21_map_block), .now(_seach_blockx_21_now));
seach_block seach_blockx_20 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_20_in_do), .start(_seach_blockx_20_start), .goal(_seach_blockx_20_goal), .data_out(_seach_blockx_20_data_out), .map_block(_seach_blockx_20_map_block), .now(_seach_blockx_20_now));
seach_block seach_blockx_19 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_19_in_do), .start(_seach_blockx_19_start), .goal(_seach_blockx_19_goal), .data_out(_seach_blockx_19_data_out), .map_block(_seach_blockx_19_map_block), .now(_seach_blockx_19_now));
seach_block seach_blockx_18 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_18_in_do), .start(_seach_blockx_18_start), .goal(_seach_blockx_18_goal), .data_out(_seach_blockx_18_data_out), .map_block(_seach_blockx_18_map_block), .now(_seach_blockx_18_now));
seach_block seach_blockx_17 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_17_in_do), .start(_seach_blockx_17_start), .goal(_seach_blockx_17_goal), .data_out(_seach_blockx_17_data_out), .map_block(_seach_blockx_17_map_block), .now(_seach_blockx_17_now));
seach_block seach_blockx_16 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_16_in_do), .start(_seach_blockx_16_start), .goal(_seach_blockx_16_goal), .data_out(_seach_blockx_16_data_out), .map_block(_seach_blockx_16_map_block), .now(_seach_blockx_16_now));
seach_block seach_blockx_15 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_15_in_do), .start(_seach_blockx_15_start), .goal(_seach_blockx_15_goal), .data_out(_seach_blockx_15_data_out), .map_block(_seach_blockx_15_map_block), .now(_seach_blockx_15_now));
seach_block seach_blockx_14 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_14_in_do), .start(_seach_blockx_14_start), .goal(_seach_blockx_14_goal), .data_out(_seach_blockx_14_data_out), .map_block(_seach_blockx_14_map_block), .now(_seach_blockx_14_now));
seach_block seach_blockx_13 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_13_in_do), .start(_seach_blockx_13_start), .goal(_seach_blockx_13_goal), .data_out(_seach_blockx_13_data_out), .map_block(_seach_blockx_13_map_block), .now(_seach_blockx_13_now));
seach_block seach_blockx_12 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_12_in_do), .start(_seach_blockx_12_start), .goal(_seach_blockx_12_goal), .data_out(_seach_blockx_12_data_out), .map_block(_seach_blockx_12_map_block), .now(_seach_blockx_12_now));
seach_block seach_blockx_11 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_11_in_do), .start(_seach_blockx_11_start), .goal(_seach_blockx_11_goal), .data_out(_seach_blockx_11_data_out), .map_block(_seach_blockx_11_map_block), .now(_seach_blockx_11_now));
seach_block seach_blockx_10 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_10_in_do), .start(_seach_blockx_10_start), .goal(_seach_blockx_10_goal), .data_out(_seach_blockx_10_data_out), .map_block(_seach_blockx_10_map_block), .now(_seach_blockx_10_now));
seach_block seach_blockx_9 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_9_in_do), .start(_seach_blockx_9_start), .goal(_seach_blockx_9_goal), .data_out(_seach_blockx_9_data_out), .map_block(_seach_blockx_9_map_block), .now(_seach_blockx_9_now));
seach_block seach_blockx_8 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_8_in_do), .start(_seach_blockx_8_start), .goal(_seach_blockx_8_goal), .data_out(_seach_blockx_8_data_out), .map_block(_seach_blockx_8_map_block), .now(_seach_blockx_8_now));
seach_block seach_blockx_7 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_7_in_do), .start(_seach_blockx_7_start), .goal(_seach_blockx_7_goal), .data_out(_seach_blockx_7_data_out), .map_block(_seach_blockx_7_map_block), .now(_seach_blockx_7_now));
seach_block seach_blockx_6 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_6_in_do), .start(_seach_blockx_6_start), .goal(_seach_blockx_6_goal), .data_out(_seach_blockx_6_data_out), .map_block(_seach_blockx_6_map_block), .now(_seach_blockx_6_now));
seach_block seach_blockx_5 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_5_in_do), .start(_seach_blockx_5_start), .goal(_seach_blockx_5_goal), .data_out(_seach_blockx_5_data_out), .map_block(_seach_blockx_5_map_block), .now(_seach_blockx_5_now));
seach_block seach_blockx_4 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_4_in_do), .start(_seach_blockx_4_start), .goal(_seach_blockx_4_goal), .data_out(_seach_blockx_4_data_out), .map_block(_seach_blockx_4_map_block), .now(_seach_blockx_4_now));
seach_block seach_blockx_3 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_3_in_do), .start(_seach_blockx_3_start), .goal(_seach_blockx_3_goal), .data_out(_seach_blockx_3_data_out), .map_block(_seach_blockx_3_map_block), .now(_seach_blockx_3_now));
seach_block seach_blockx_2 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_2_in_do), .start(_seach_blockx_2_start), .goal(_seach_blockx_2_goal), .data_out(_seach_blockx_2_data_out), .map_block(_seach_blockx_2_map_block), .now(_seach_blockx_2_now));
seach_block seach_blockx_1 (.m_clock(m_clock), .p_reset( p_reset), .in_do(_seach_blockx_1_in_do), .start(_seach_blockx_1_start), .goal(_seach_blockx_1_goal), .data_out(_seach_blockx_1_data_out), .map_block(_seach_blockx_1_map_block), .now(_seach_blockx_1_now));

   assign  _seach_blockx_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in17:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00010001:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_in_do)
  begin
#1 if (_seach_blockx_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 14 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_in_do = (in_do|_reg_1);
   assign  _seach_blockx_p_reset = p_reset;
   assign  _seach_blockx_m_clock = m_clock;
   assign  _seach_blockx_195_in_do = 1'b0;
   assign  _seach_blockx_195_p_reset = p_reset;
   assign  _seach_blockx_195_m_clock = m_clock;
   assign  _seach_blockx_194_in_do = 1'b0;
   assign  _seach_blockx_194_p_reset = p_reset;
   assign  _seach_blockx_194_m_clock = m_clock;
   assign  _seach_blockx_193_in_do = 1'b0;
   assign  _seach_blockx_193_p_reset = p_reset;
   assign  _seach_blockx_193_m_clock = m_clock;
   assign  _seach_blockx_192_in_do = 1'b0;
   assign  _seach_blockx_192_p_reset = p_reset;
   assign  _seach_blockx_192_m_clock = m_clock;
   assign  _seach_blockx_191_in_do = 1'b0;
   assign  _seach_blockx_191_p_reset = p_reset;
   assign  _seach_blockx_191_m_clock = m_clock;
   assign  _seach_blockx_190_in_do = 1'b0;
   assign  _seach_blockx_190_p_reset = p_reset;
   assign  _seach_blockx_190_m_clock = m_clock;
   assign  _seach_blockx_189_in_do = 1'b0;
   assign  _seach_blockx_189_p_reset = p_reset;
   assign  _seach_blockx_189_m_clock = m_clock;
   assign  _seach_blockx_188_in_do = 1'b0;
   assign  _seach_blockx_188_p_reset = p_reset;
   assign  _seach_blockx_188_m_clock = m_clock;
   assign  _seach_blockx_187_in_do = 1'b0;
   assign  _seach_blockx_187_p_reset = p_reset;
   assign  _seach_blockx_187_m_clock = m_clock;
   assign  _seach_blockx_186_in_do = 1'b0;
   assign  _seach_blockx_186_p_reset = p_reset;
   assign  _seach_blockx_186_m_clock = m_clock;
   assign  _seach_blockx_185_in_do = 1'b0;
   assign  _seach_blockx_185_p_reset = p_reset;
   assign  _seach_blockx_185_m_clock = m_clock;
   assign  _seach_blockx_184_in_do = 1'b0;
   assign  _seach_blockx_184_p_reset = p_reset;
   assign  _seach_blockx_184_m_clock = m_clock;
   assign  _seach_blockx_183_in_do = 1'b0;
   assign  _seach_blockx_183_p_reset = p_reset;
   assign  _seach_blockx_183_m_clock = m_clock;
   assign  _seach_blockx_182_in_do = 1'b0;
   assign  _seach_blockx_182_p_reset = p_reset;
   assign  _seach_blockx_182_m_clock = m_clock;
   assign  _seach_blockx_181_in_do = 1'b0;
   assign  _seach_blockx_181_p_reset = p_reset;
   assign  _seach_blockx_181_m_clock = m_clock;
   assign  _seach_blockx_180_in_do = 1'b0;
   assign  _seach_blockx_180_p_reset = p_reset;
   assign  _seach_blockx_180_m_clock = m_clock;
   assign  _seach_blockx_179_in_do = 1'b0;
   assign  _seach_blockx_179_p_reset = p_reset;
   assign  _seach_blockx_179_m_clock = m_clock;
   assign  _seach_blockx_178_in_do = 1'b0;
   assign  _seach_blockx_178_p_reset = p_reset;
   assign  _seach_blockx_178_m_clock = m_clock;
   assign  _seach_blockx_177_in_do = 1'b0;
   assign  _seach_blockx_177_p_reset = p_reset;
   assign  _seach_blockx_177_m_clock = m_clock;
   assign  _seach_blockx_176_in_do = 1'b0;
   assign  _seach_blockx_176_p_reset = p_reset;
   assign  _seach_blockx_176_m_clock = m_clock;
   assign  _seach_blockx_175_in_do = 1'b0;
   assign  _seach_blockx_175_p_reset = p_reset;
   assign  _seach_blockx_175_m_clock = m_clock;
   assign  _seach_blockx_174_in_do = 1'b0;
   assign  _seach_blockx_174_p_reset = p_reset;
   assign  _seach_blockx_174_m_clock = m_clock;
   assign  _seach_blockx_173_in_do = 1'b0;
   assign  _seach_blockx_173_p_reset = p_reset;
   assign  _seach_blockx_173_m_clock = m_clock;
   assign  _seach_blockx_172_in_do = 1'b0;
   assign  _seach_blockx_172_p_reset = p_reset;
   assign  _seach_blockx_172_m_clock = m_clock;
   assign  _seach_blockx_171_in_do = 1'b0;
   assign  _seach_blockx_171_p_reset = p_reset;
   assign  _seach_blockx_171_m_clock = m_clock;
   assign  _seach_blockx_170_in_do = 1'b0;
   assign  _seach_blockx_170_p_reset = p_reset;
   assign  _seach_blockx_170_m_clock = m_clock;
   assign  _seach_blockx_169_in_do = 1'b0;
   assign  _seach_blockx_169_p_reset = p_reset;
   assign  _seach_blockx_169_m_clock = m_clock;
   assign  _seach_blockx_168_in_do = 1'b0;
   assign  _seach_blockx_168_p_reset = p_reset;
   assign  _seach_blockx_168_m_clock = m_clock;
   assign  _seach_blockx_167_in_do = 1'b0;
   assign  _seach_blockx_167_p_reset = p_reset;
   assign  _seach_blockx_167_m_clock = m_clock;
   assign  _seach_blockx_166_in_do = 1'b0;
   assign  _seach_blockx_166_p_reset = p_reset;
   assign  _seach_blockx_166_m_clock = m_clock;
   assign  _seach_blockx_165_in_do = 1'b0;
   assign  _seach_blockx_165_p_reset = p_reset;
   assign  _seach_blockx_165_m_clock = m_clock;
   assign  _seach_blockx_164_in_do = 1'b0;
   assign  _seach_blockx_164_p_reset = p_reset;
   assign  _seach_blockx_164_m_clock = m_clock;
   assign  _seach_blockx_163_in_do = 1'b0;
   assign  _seach_blockx_163_p_reset = p_reset;
   assign  _seach_blockx_163_m_clock = m_clock;
   assign  _seach_blockx_162_in_do = 1'b0;
   assign  _seach_blockx_162_p_reset = p_reset;
   assign  _seach_blockx_162_m_clock = m_clock;
   assign  _seach_blockx_161_in_do = 1'b0;
   assign  _seach_blockx_161_p_reset = p_reset;
   assign  _seach_blockx_161_m_clock = m_clock;
   assign  _seach_blockx_160_in_do = 1'b0;
   assign  _seach_blockx_160_p_reset = p_reset;
   assign  _seach_blockx_160_m_clock = m_clock;
   assign  _seach_blockx_159_in_do = 1'b0;
   assign  _seach_blockx_159_p_reset = p_reset;
   assign  _seach_blockx_159_m_clock = m_clock;
   assign  _seach_blockx_158_in_do = 1'b0;
   assign  _seach_blockx_158_p_reset = p_reset;
   assign  _seach_blockx_158_m_clock = m_clock;
   assign  _seach_blockx_157_in_do = 1'b0;
   assign  _seach_blockx_157_p_reset = p_reset;
   assign  _seach_blockx_157_m_clock = m_clock;
   assign  _seach_blockx_156_in_do = 1'b0;
   assign  _seach_blockx_156_p_reset = p_reset;
   assign  _seach_blockx_156_m_clock = m_clock;
   assign  _seach_blockx_155_in_do = 1'b0;
   assign  _seach_blockx_155_p_reset = p_reset;
   assign  _seach_blockx_155_m_clock = m_clock;
   assign  _seach_blockx_154_in_do = 1'b0;
   assign  _seach_blockx_154_p_reset = p_reset;
   assign  _seach_blockx_154_m_clock = m_clock;
   assign  _seach_blockx_153_in_do = 1'b0;
   assign  _seach_blockx_153_p_reset = p_reset;
   assign  _seach_blockx_153_m_clock = m_clock;
   assign  _seach_blockx_152_in_do = 1'b0;
   assign  _seach_blockx_152_p_reset = p_reset;
   assign  _seach_blockx_152_m_clock = m_clock;
   assign  _seach_blockx_151_in_do = 1'b0;
   assign  _seach_blockx_151_p_reset = p_reset;
   assign  _seach_blockx_151_m_clock = m_clock;
   assign  _seach_blockx_150_in_do = 1'b0;
   assign  _seach_blockx_150_p_reset = p_reset;
   assign  _seach_blockx_150_m_clock = m_clock;
   assign  _seach_blockx_149_in_do = 1'b0;
   assign  _seach_blockx_149_p_reset = p_reset;
   assign  _seach_blockx_149_m_clock = m_clock;
   assign  _seach_blockx_148_in_do = 1'b0;
   assign  _seach_blockx_148_p_reset = p_reset;
   assign  _seach_blockx_148_m_clock = m_clock;
   assign  _seach_blockx_147_in_do = 1'b0;
   assign  _seach_blockx_147_p_reset = p_reset;
   assign  _seach_blockx_147_m_clock = m_clock;
   assign  _seach_blockx_146_in_do = 1'b0;
   assign  _seach_blockx_146_p_reset = p_reset;
   assign  _seach_blockx_146_m_clock = m_clock;
   assign  _seach_blockx_145_in_do = 1'b0;
   assign  _seach_blockx_145_p_reset = p_reset;
   assign  _seach_blockx_145_m_clock = m_clock;
   assign  _seach_blockx_144_in_do = 1'b0;
   assign  _seach_blockx_144_p_reset = p_reset;
   assign  _seach_blockx_144_m_clock = m_clock;
   assign  _seach_blockx_143_in_do = 1'b0;
   assign  _seach_blockx_143_p_reset = p_reset;
   assign  _seach_blockx_143_m_clock = m_clock;
   assign  _seach_blockx_142_in_do = 1'b0;
   assign  _seach_blockx_142_p_reset = p_reset;
   assign  _seach_blockx_142_m_clock = m_clock;
   assign  _seach_blockx_141_in_do = 1'b0;
   assign  _seach_blockx_141_p_reset = p_reset;
   assign  _seach_blockx_141_m_clock = m_clock;
   assign  _seach_blockx_140_in_do = 1'b0;
   assign  _seach_blockx_140_p_reset = p_reset;
   assign  _seach_blockx_140_m_clock = m_clock;
   assign  _seach_blockx_139_in_do = 1'b0;
   assign  _seach_blockx_139_p_reset = p_reset;
   assign  _seach_blockx_139_m_clock = m_clock;
   assign  _seach_blockx_138_in_do = 1'b0;
   assign  _seach_blockx_138_p_reset = p_reset;
   assign  _seach_blockx_138_m_clock = m_clock;
   assign  _seach_blockx_137_in_do = 1'b0;
   assign  _seach_blockx_137_p_reset = p_reset;
   assign  _seach_blockx_137_m_clock = m_clock;
   assign  _seach_blockx_136_in_do = 1'b0;
   assign  _seach_blockx_136_p_reset = p_reset;
   assign  _seach_blockx_136_m_clock = m_clock;
   assign  _seach_blockx_135_in_do = 1'b0;
   assign  _seach_blockx_135_p_reset = p_reset;
   assign  _seach_blockx_135_m_clock = m_clock;
   assign  _seach_blockx_134_in_do = 1'b0;
   assign  _seach_blockx_134_p_reset = p_reset;
   assign  _seach_blockx_134_m_clock = m_clock;
   assign  _seach_blockx_133_in_do = 1'b0;
   assign  _seach_blockx_133_p_reset = p_reset;
   assign  _seach_blockx_133_m_clock = m_clock;
   assign  _seach_blockx_132_in_do = 1'b0;
   assign  _seach_blockx_132_p_reset = p_reset;
   assign  _seach_blockx_132_m_clock = m_clock;
   assign  _seach_blockx_131_in_do = 1'b0;
   assign  _seach_blockx_131_p_reset = p_reset;
   assign  _seach_blockx_131_m_clock = m_clock;
   assign  _seach_blockx_130_in_do = 1'b0;
   assign  _seach_blockx_130_p_reset = p_reset;
   assign  _seach_blockx_130_m_clock = m_clock;
   assign  _seach_blockx_129_in_do = 1'b0;
   assign  _seach_blockx_129_p_reset = p_reset;
   assign  _seach_blockx_129_m_clock = m_clock;
   assign  _seach_blockx_128_in_do = 1'b0;
   assign  _seach_blockx_128_p_reset = p_reset;
   assign  _seach_blockx_128_m_clock = m_clock;
   assign  _seach_blockx_127_in_do = 1'b0;
   assign  _seach_blockx_127_p_reset = p_reset;
   assign  _seach_blockx_127_m_clock = m_clock;
   assign  _seach_blockx_126_in_do = 1'b0;
   assign  _seach_blockx_126_p_reset = p_reset;
   assign  _seach_blockx_126_m_clock = m_clock;
   assign  _seach_blockx_125_in_do = 1'b0;
   assign  _seach_blockx_125_p_reset = p_reset;
   assign  _seach_blockx_125_m_clock = m_clock;
   assign  _seach_blockx_124_in_do = 1'b0;
   assign  _seach_blockx_124_p_reset = p_reset;
   assign  _seach_blockx_124_m_clock = m_clock;
   assign  _seach_blockx_123_in_do = 1'b0;
   assign  _seach_blockx_123_p_reset = p_reset;
   assign  _seach_blockx_123_m_clock = m_clock;
   assign  _seach_blockx_122_in_do = 1'b0;
   assign  _seach_blockx_122_p_reset = p_reset;
   assign  _seach_blockx_122_m_clock = m_clock;
   assign  _seach_blockx_121_in_do = 1'b0;
   assign  _seach_blockx_121_p_reset = p_reset;
   assign  _seach_blockx_121_m_clock = m_clock;
   assign  _seach_blockx_120_in_do = 1'b0;
   assign  _seach_blockx_120_p_reset = p_reset;
   assign  _seach_blockx_120_m_clock = m_clock;
   assign  _seach_blockx_119_in_do = 1'b0;
   assign  _seach_blockx_119_p_reset = p_reset;
   assign  _seach_blockx_119_m_clock = m_clock;
   assign  _seach_blockx_118_in_do = 1'b0;
   assign  _seach_blockx_118_p_reset = p_reset;
   assign  _seach_blockx_118_m_clock = m_clock;
   assign  _seach_blockx_117_in_do = 1'b0;
   assign  _seach_blockx_117_p_reset = p_reset;
   assign  _seach_blockx_117_m_clock = m_clock;
   assign  _seach_blockx_116_in_do = 1'b0;
   assign  _seach_blockx_116_p_reset = p_reset;
   assign  _seach_blockx_116_m_clock = m_clock;
   assign  _seach_blockx_115_in_do = 1'b0;
   assign  _seach_blockx_115_p_reset = p_reset;
   assign  _seach_blockx_115_m_clock = m_clock;
   assign  _seach_blockx_114_in_do = 1'b0;
   assign  _seach_blockx_114_p_reset = p_reset;
   assign  _seach_blockx_114_m_clock = m_clock;
   assign  _seach_blockx_113_in_do = 1'b0;
   assign  _seach_blockx_113_p_reset = p_reset;
   assign  _seach_blockx_113_m_clock = m_clock;
   assign  _seach_blockx_112_in_do = 1'b0;
   assign  _seach_blockx_112_p_reset = p_reset;
   assign  _seach_blockx_112_m_clock = m_clock;
   assign  _seach_blockx_111_in_do = 1'b0;
   assign  _seach_blockx_111_p_reset = p_reset;
   assign  _seach_blockx_111_m_clock = m_clock;
   assign  _seach_blockx_110_in_do = 1'b0;
   assign  _seach_blockx_110_p_reset = p_reset;
   assign  _seach_blockx_110_m_clock = m_clock;
   assign  _seach_blockx_109_in_do = 1'b0;
   assign  _seach_blockx_109_p_reset = p_reset;
   assign  _seach_blockx_109_m_clock = m_clock;
   assign  _seach_blockx_108_in_do = 1'b0;
   assign  _seach_blockx_108_p_reset = p_reset;
   assign  _seach_blockx_108_m_clock = m_clock;
   assign  _seach_blockx_107_in_do = 1'b0;
   assign  _seach_blockx_107_p_reset = p_reset;
   assign  _seach_blockx_107_m_clock = m_clock;
   assign  _seach_blockx_106_in_do = 1'b0;
   assign  _seach_blockx_106_p_reset = p_reset;
   assign  _seach_blockx_106_m_clock = m_clock;
   assign  _seach_blockx_105_in_do = 1'b0;
   assign  _seach_blockx_105_p_reset = p_reset;
   assign  _seach_blockx_105_m_clock = m_clock;
   assign  _seach_blockx_104_in_do = 1'b0;
   assign  _seach_blockx_104_p_reset = p_reset;
   assign  _seach_blockx_104_m_clock = m_clock;
   assign  _seach_blockx_103_in_do = 1'b0;
   assign  _seach_blockx_103_p_reset = p_reset;
   assign  _seach_blockx_103_m_clock = m_clock;
   assign  _seach_blockx_102_in_do = 1'b0;
   assign  _seach_blockx_102_p_reset = p_reset;
   assign  _seach_blockx_102_m_clock = m_clock;
   assign  _seach_blockx_101_in_do = 1'b0;
   assign  _seach_blockx_101_p_reset = p_reset;
   assign  _seach_blockx_101_m_clock = m_clock;
   assign  _seach_blockx_100_in_do = 1'b0;
   assign  _seach_blockx_100_p_reset = p_reset;
   assign  _seach_blockx_100_m_clock = m_clock;
   assign  _seach_blockx_99_in_do = 1'b0;
   assign  _seach_blockx_99_p_reset = p_reset;
   assign  _seach_blockx_99_m_clock = m_clock;
   assign  _seach_blockx_98_in_do = 1'b0;
   assign  _seach_blockx_98_p_reset = p_reset;
   assign  _seach_blockx_98_m_clock = m_clock;
   assign  _seach_blockx_97_in_do = 1'b0;
   assign  _seach_blockx_97_p_reset = p_reset;
   assign  _seach_blockx_97_m_clock = m_clock;
   assign  _seach_blockx_96_in_do = 1'b0;
   assign  _seach_blockx_96_p_reset = p_reset;
   assign  _seach_blockx_96_m_clock = m_clock;
   assign  _seach_blockx_95_in_do = 1'b0;
   assign  _seach_blockx_95_p_reset = p_reset;
   assign  _seach_blockx_95_m_clock = m_clock;
   assign  _seach_blockx_94_in_do = 1'b0;
   assign  _seach_blockx_94_p_reset = p_reset;
   assign  _seach_blockx_94_m_clock = m_clock;
   assign  _seach_blockx_93_in_do = 1'b0;
   assign  _seach_blockx_93_p_reset = p_reset;
   assign  _seach_blockx_93_m_clock = m_clock;
   assign  _seach_blockx_92_in_do = 1'b0;
   assign  _seach_blockx_92_p_reset = p_reset;
   assign  _seach_blockx_92_m_clock = m_clock;
   assign  _seach_blockx_91_in_do = 1'b0;
   assign  _seach_blockx_91_p_reset = p_reset;
   assign  _seach_blockx_91_m_clock = m_clock;
   assign  _seach_blockx_90_in_do = 1'b0;
   assign  _seach_blockx_90_p_reset = p_reset;
   assign  _seach_blockx_90_m_clock = m_clock;
   assign  _seach_blockx_89_in_do = 1'b0;
   assign  _seach_blockx_89_p_reset = p_reset;
   assign  _seach_blockx_89_m_clock = m_clock;
   assign  _seach_blockx_88_in_do = 1'b0;
   assign  _seach_blockx_88_p_reset = p_reset;
   assign  _seach_blockx_88_m_clock = m_clock;
   assign  _seach_blockx_87_in_do = 1'b0;
   assign  _seach_blockx_87_p_reset = p_reset;
   assign  _seach_blockx_87_m_clock = m_clock;
   assign  _seach_blockx_86_in_do = 1'b0;
   assign  _seach_blockx_86_p_reset = p_reset;
   assign  _seach_blockx_86_m_clock = m_clock;
   assign  _seach_blockx_85_in_do = 1'b0;
   assign  _seach_blockx_85_p_reset = p_reset;
   assign  _seach_blockx_85_m_clock = m_clock;
   assign  _seach_blockx_84_in_do = 1'b0;
   assign  _seach_blockx_84_p_reset = p_reset;
   assign  _seach_blockx_84_m_clock = m_clock;
   assign  _seach_blockx_83_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in110:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_83_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01101110:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_83_in_do)
  begin
#1 if (_seach_blockx_83_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_83_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 97 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_83_in_do = (in_do|_reg_1);
   assign  _seach_blockx_83_p_reset = p_reset;
   assign  _seach_blockx_83_m_clock = m_clock;
   assign  _seach_blockx_82_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in109:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_82_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01101101:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_82_in_do)
  begin
#1 if (_seach_blockx_82_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_82_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 96 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_82_in_do = (in_do|_reg_1);
   assign  _seach_blockx_82_p_reset = p_reset;
   assign  _seach_blockx_82_m_clock = m_clock;
   assign  _seach_blockx_81_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in108:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_81_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01101100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_81_in_do)
  begin
#1 if (_seach_blockx_81_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_81_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 95 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_81_in_do = (in_do|_reg_1);
   assign  _seach_blockx_81_p_reset = p_reset;
   assign  _seach_blockx_81_m_clock = m_clock;
   assign  _seach_blockx_80_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in107:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_80_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01101011:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_80_in_do)
  begin
#1 if (_seach_blockx_80_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_80_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 94 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_80_in_do = (in_do|_reg_1);
   assign  _seach_blockx_80_p_reset = p_reset;
   assign  _seach_blockx_80_m_clock = m_clock;
   assign  _seach_blockx_79_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in106:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_79_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01101010:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_79_in_do)
  begin
#1 if (_seach_blockx_79_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_79_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 93 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_79_in_do = (in_do|_reg_1);
   assign  _seach_blockx_79_p_reset = p_reset;
   assign  _seach_blockx_79_m_clock = m_clock;
   assign  _seach_blockx_78_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in105:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_78_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01101001:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_78_in_do)
  begin
#1 if (_seach_blockx_78_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_78_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 92 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_78_in_do = (in_do|_reg_1);
   assign  _seach_blockx_78_p_reset = p_reset;
   assign  _seach_blockx_78_m_clock = m_clock;
   assign  _seach_blockx_77_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in104:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_77_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01101000:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_77_in_do)
  begin
#1 if (_seach_blockx_77_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_77_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 91 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_77_in_do = (in_do|_reg_1);
   assign  _seach_blockx_77_p_reset = p_reset;
   assign  _seach_blockx_77_m_clock = m_clock;
   assign  _seach_blockx_76_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in103:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_76_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01100111:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_76_in_do)
  begin
#1 if (_seach_blockx_76_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_76_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 90 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_76_in_do = (in_do|_reg_1);
   assign  _seach_blockx_76_p_reset = p_reset;
   assign  _seach_blockx_76_m_clock = m_clock;
   assign  _seach_blockx_75_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in102:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_75_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01100110:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_75_in_do)
  begin
#1 if (_seach_blockx_75_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_75_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 89 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_75_in_do = (in_do|_reg_1);
   assign  _seach_blockx_75_p_reset = p_reset;
   assign  _seach_blockx_75_m_clock = m_clock;
   assign  _seach_blockx_74_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in101:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_74_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01100101:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_74_in_do)
  begin
#1 if (_seach_blockx_74_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_74_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 88 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_74_in_do = (in_do|_reg_1);
   assign  _seach_blockx_74_p_reset = p_reset;
   assign  _seach_blockx_74_m_clock = m_clock;
   assign  _seach_blockx_73_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_73_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01100100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_73_in_do)
  begin
#1 if (_seach_blockx_73_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_73_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 87 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_73_in_do = (in_do|_reg_1);
   assign  _seach_blockx_73_p_reset = p_reset;
   assign  _seach_blockx_73_m_clock = m_clock;
   assign  _seach_blockx_72_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in99:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_72_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01100011:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_72_in_do)
  begin
#1 if (_seach_blockx_72_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_72_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 86 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_72_in_do = (in_do|_reg_1);
   assign  _seach_blockx_72_p_reset = p_reset;
   assign  _seach_blockx_72_m_clock = m_clock;
   assign  _seach_blockx_71_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in98:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_71_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01100010:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_71_in_do)
  begin
#1 if (_seach_blockx_71_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_71_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 85 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_71_in_do = (in_do|_reg_1);
   assign  _seach_blockx_71_p_reset = p_reset;
   assign  _seach_blockx_71_m_clock = m_clock;
   assign  _seach_blockx_70_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in97:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_70_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01100001:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_70_in_do)
  begin
#1 if (_seach_blockx_70_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_70_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 84 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_70_in_do = (in_do|_reg_1);
   assign  _seach_blockx_70_p_reset = p_reset;
   assign  _seach_blockx_70_m_clock = m_clock;
   assign  _seach_blockx_69_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in94:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_69_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01011110:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_69_in_do)
  begin
#1 if (_seach_blockx_69_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_69_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 83 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_69_in_do = (in_do|_reg_1);
   assign  _seach_blockx_69_p_reset = p_reset;
   assign  _seach_blockx_69_m_clock = m_clock;
   assign  _seach_blockx_68_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in93:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_68_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01011101:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_68_in_do)
  begin
#1 if (_seach_blockx_68_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_68_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 82 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_68_in_do = (in_do|_reg_1);
   assign  _seach_blockx_68_p_reset = p_reset;
   assign  _seach_blockx_68_m_clock = m_clock;
   assign  _seach_blockx_67_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in92:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_67_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01011100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_67_in_do)
  begin
#1 if (_seach_blockx_67_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_67_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 81 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_67_in_do = (in_do|_reg_1);
   assign  _seach_blockx_67_p_reset = p_reset;
   assign  _seach_blockx_67_m_clock = m_clock;
   assign  _seach_blockx_66_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in91:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_66_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01011011:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_66_in_do)
  begin
#1 if (_seach_blockx_66_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_66_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 80 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_66_in_do = (in_do|_reg_1);
   assign  _seach_blockx_66_p_reset = p_reset;
   assign  _seach_blockx_66_m_clock = m_clock;
   assign  _seach_blockx_65_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in90:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_65_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01011010:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_65_in_do)
  begin
#1 if (_seach_blockx_65_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_65_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 79 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_65_in_do = (in_do|_reg_1);
   assign  _seach_blockx_65_p_reset = p_reset;
   assign  _seach_blockx_65_m_clock = m_clock;
   assign  _seach_blockx_64_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in89:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_64_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01011001:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_64_in_do)
  begin
#1 if (_seach_blockx_64_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_64_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 78 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_64_in_do = (in_do|_reg_1);
   assign  _seach_blockx_64_p_reset = p_reset;
   assign  _seach_blockx_64_m_clock = m_clock;
   assign  _seach_blockx_63_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in88:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_63_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01011000:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_63_in_do)
  begin
#1 if (_seach_blockx_63_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_63_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 77 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_63_in_do = (in_do|_reg_1);
   assign  _seach_blockx_63_p_reset = p_reset;
   assign  _seach_blockx_63_m_clock = m_clock;
   assign  _seach_blockx_62_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in87:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_62_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01010111:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_62_in_do)
  begin
#1 if (_seach_blockx_62_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_62_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 76 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_62_in_do = (in_do|_reg_1);
   assign  _seach_blockx_62_p_reset = p_reset;
   assign  _seach_blockx_62_m_clock = m_clock;
   assign  _seach_blockx_61_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in86:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_61_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01010110:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_61_in_do)
  begin
#1 if (_seach_blockx_61_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_61_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 75 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_61_in_do = (in_do|_reg_1);
   assign  _seach_blockx_61_p_reset = p_reset;
   assign  _seach_blockx_61_m_clock = m_clock;
   assign  _seach_blockx_60_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in85:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_60_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01010101:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_60_in_do)
  begin
#1 if (_seach_blockx_60_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_60_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 74 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_60_in_do = (in_do|_reg_1);
   assign  _seach_blockx_60_p_reset = p_reset;
   assign  _seach_blockx_60_m_clock = m_clock;
   assign  _seach_blockx_59_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in84:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_59_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01010100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_59_in_do)
  begin
#1 if (_seach_blockx_59_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_59_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 73 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_59_in_do = (in_do|_reg_1);
   assign  _seach_blockx_59_p_reset = p_reset;
   assign  _seach_blockx_59_m_clock = m_clock;
   assign  _seach_blockx_58_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in83:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_58_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01010011:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_58_in_do)
  begin
#1 if (_seach_blockx_58_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_58_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 72 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_58_in_do = (in_do|_reg_1);
   assign  _seach_blockx_58_p_reset = p_reset;
   assign  _seach_blockx_58_m_clock = m_clock;
   assign  _seach_blockx_57_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in82:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_57_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01010010:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_57_in_do)
  begin
#1 if (_seach_blockx_57_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_57_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 71 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_57_in_do = (in_do|_reg_1);
   assign  _seach_blockx_57_p_reset = p_reset;
   assign  _seach_blockx_57_m_clock = m_clock;
   assign  _seach_blockx_56_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in81:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_56_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01010001:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_56_in_do)
  begin
#1 if (_seach_blockx_56_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_56_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 70 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_56_in_do = (in_do|_reg_1);
   assign  _seach_blockx_56_p_reset = p_reset;
   assign  _seach_blockx_56_m_clock = m_clock;
   assign  _seach_blockx_55_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in78:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_55_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01001110:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_55_in_do)
  begin
#1 if (_seach_blockx_55_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_55_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 69 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_55_in_do = (in_do|_reg_1);
   assign  _seach_blockx_55_p_reset = p_reset;
   assign  _seach_blockx_55_m_clock = m_clock;
   assign  _seach_blockx_54_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in77:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_54_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01001101:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_54_in_do)
  begin
#1 if (_seach_blockx_54_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_54_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 68 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_54_in_do = (in_do|_reg_1);
   assign  _seach_blockx_54_p_reset = p_reset;
   assign  _seach_blockx_54_m_clock = m_clock;
   assign  _seach_blockx_53_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in76:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_53_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01001100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_53_in_do)
  begin
#1 if (_seach_blockx_53_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_53_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 67 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_53_in_do = (in_do|_reg_1);
   assign  _seach_blockx_53_p_reset = p_reset;
   assign  _seach_blockx_53_m_clock = m_clock;
   assign  _seach_blockx_52_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in75:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_52_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01001011:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_52_in_do)
  begin
#1 if (_seach_blockx_52_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_52_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 66 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_52_in_do = (in_do|_reg_1);
   assign  _seach_blockx_52_p_reset = p_reset;
   assign  _seach_blockx_52_m_clock = m_clock;
   assign  _seach_blockx_51_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in74:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_51_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01001010:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_51_in_do)
  begin
#1 if (_seach_blockx_51_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_51_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 65 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_51_in_do = (in_do|_reg_1);
   assign  _seach_blockx_51_p_reset = p_reset;
   assign  _seach_blockx_51_m_clock = m_clock;
   assign  _seach_blockx_50_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in73:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_50_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01001001:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_50_in_do)
  begin
#1 if (_seach_blockx_50_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_50_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 64 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_50_in_do = (in_do|_reg_1);
   assign  _seach_blockx_50_p_reset = p_reset;
   assign  _seach_blockx_50_m_clock = m_clock;
   assign  _seach_blockx_49_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in72:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_49_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01001000:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_49_in_do)
  begin
#1 if (_seach_blockx_49_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_49_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 63 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_49_in_do = (in_do|_reg_1);
   assign  _seach_blockx_49_p_reset = p_reset;
   assign  _seach_blockx_49_m_clock = m_clock;
   assign  _seach_blockx_48_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in71:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_48_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01000111:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_48_in_do)
  begin
#1 if (_seach_blockx_48_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_48_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 62 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_48_in_do = (in_do|_reg_1);
   assign  _seach_blockx_48_p_reset = p_reset;
   assign  _seach_blockx_48_m_clock = m_clock;
   assign  _seach_blockx_47_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in70:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_47_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01000110:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_47_in_do)
  begin
#1 if (_seach_blockx_47_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_47_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 61 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_47_in_do = (in_do|_reg_1);
   assign  _seach_blockx_47_p_reset = p_reset;
   assign  _seach_blockx_47_m_clock = m_clock;
   assign  _seach_blockx_46_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in69:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_46_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01000101:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_46_in_do)
  begin
#1 if (_seach_blockx_46_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_46_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 60 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_46_in_do = (in_do|_reg_1);
   assign  _seach_blockx_46_p_reset = p_reset;
   assign  _seach_blockx_46_m_clock = m_clock;
   assign  _seach_blockx_45_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in68:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_45_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01000100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_45_in_do)
  begin
#1 if (_seach_blockx_45_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_45_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 59 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_45_in_do = (in_do|_reg_1);
   assign  _seach_blockx_45_p_reset = p_reset;
   assign  _seach_blockx_45_m_clock = m_clock;
   assign  _seach_blockx_44_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in67:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_44_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01000011:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_44_in_do)
  begin
#1 if (_seach_blockx_44_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_44_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 58 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_44_in_do = (in_do|_reg_1);
   assign  _seach_blockx_44_p_reset = p_reset;
   assign  _seach_blockx_44_m_clock = m_clock;
   assign  _seach_blockx_43_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in66:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_43_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01000010:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_43_in_do)
  begin
#1 if (_seach_blockx_43_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_43_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 57 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_43_in_do = (in_do|_reg_1);
   assign  _seach_blockx_43_p_reset = p_reset;
   assign  _seach_blockx_43_m_clock = m_clock;
   assign  _seach_blockx_42_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in65:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_42_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b01000001:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_42_in_do)
  begin
#1 if (_seach_blockx_42_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_42_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 56 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_42_in_do = (in_do|_reg_1);
   assign  _seach_blockx_42_p_reset = p_reset;
   assign  _seach_blockx_42_m_clock = m_clock;
   assign  _seach_blockx_41_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in62:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_41_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00111110:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_41_in_do)
  begin
#1 if (_seach_blockx_41_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_41_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 55 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_41_in_do = (in_do|_reg_1);
   assign  _seach_blockx_41_p_reset = p_reset;
   assign  _seach_blockx_41_m_clock = m_clock;
   assign  _seach_blockx_40_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in61:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_40_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00111101:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_40_in_do)
  begin
#1 if (_seach_blockx_40_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_40_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 54 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_40_in_do = (in_do|_reg_1);
   assign  _seach_blockx_40_p_reset = p_reset;
   assign  _seach_blockx_40_m_clock = m_clock;
   assign  _seach_blockx_39_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in60:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_39_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00111100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_39_in_do)
  begin
#1 if (_seach_blockx_39_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_39_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 53 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_39_in_do = (in_do|_reg_1);
   assign  _seach_blockx_39_p_reset = p_reset;
   assign  _seach_blockx_39_m_clock = m_clock;
   assign  _seach_blockx_38_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in59:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_38_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00111011:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_38_in_do)
  begin
#1 if (_seach_blockx_38_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_38_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 52 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_38_in_do = (in_do|_reg_1);
   assign  _seach_blockx_38_p_reset = p_reset;
   assign  _seach_blockx_38_m_clock = m_clock;
   assign  _seach_blockx_37_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in58:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_37_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00111010:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_37_in_do)
  begin
#1 if (_seach_blockx_37_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_37_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 51 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_37_in_do = (in_do|_reg_1);
   assign  _seach_blockx_37_p_reset = p_reset;
   assign  _seach_blockx_37_m_clock = m_clock;
   assign  _seach_blockx_36_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in57:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_36_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00111001:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_36_in_do)
  begin
#1 if (_seach_blockx_36_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_36_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 50 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_36_in_do = (in_do|_reg_1);
   assign  _seach_blockx_36_p_reset = p_reset;
   assign  _seach_blockx_36_m_clock = m_clock;
   assign  _seach_blockx_35_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in56:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_35_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00111000:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_35_in_do)
  begin
#1 if (_seach_blockx_35_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_35_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 49 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_35_in_do = (in_do|_reg_1);
   assign  _seach_blockx_35_p_reset = p_reset;
   assign  _seach_blockx_35_m_clock = m_clock;
   assign  _seach_blockx_34_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in55:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_34_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00110111:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_34_in_do)
  begin
#1 if (_seach_blockx_34_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_34_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 48 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_34_in_do = (in_do|_reg_1);
   assign  _seach_blockx_34_p_reset = p_reset;
   assign  _seach_blockx_34_m_clock = m_clock;
   assign  _seach_blockx_33_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in54:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_33_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00110110:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_33_in_do)
  begin
#1 if (_seach_blockx_33_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_33_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 47 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_33_in_do = (in_do|_reg_1);
   assign  _seach_blockx_33_p_reset = p_reset;
   assign  _seach_blockx_33_m_clock = m_clock;
   assign  _seach_blockx_32_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in53:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_32_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00110101:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_32_in_do)
  begin
#1 if (_seach_blockx_32_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_32_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 46 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_32_in_do = (in_do|_reg_1);
   assign  _seach_blockx_32_p_reset = p_reset;
   assign  _seach_blockx_32_m_clock = m_clock;
   assign  _seach_blockx_31_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in52:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_31_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00110100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_31_in_do)
  begin
#1 if (_seach_blockx_31_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_31_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 45 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_31_in_do = (in_do|_reg_1);
   assign  _seach_blockx_31_p_reset = p_reset;
   assign  _seach_blockx_31_m_clock = m_clock;
   assign  _seach_blockx_30_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in51:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_30_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00110011:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_30_in_do)
  begin
#1 if (_seach_blockx_30_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_30_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 44 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_30_in_do = (in_do|_reg_1);
   assign  _seach_blockx_30_p_reset = p_reset;
   assign  _seach_blockx_30_m_clock = m_clock;
   assign  _seach_blockx_29_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in50:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_29_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00110010:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_29_in_do)
  begin
#1 if (_seach_blockx_29_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_29_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 43 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_29_in_do = (in_do|_reg_1);
   assign  _seach_blockx_29_p_reset = p_reset;
   assign  _seach_blockx_29_m_clock = m_clock;
   assign  _seach_blockx_28_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in49:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_28_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00110001:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_28_in_do)
  begin
#1 if (_seach_blockx_28_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_28_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 42 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_28_in_do = (in_do|_reg_1);
   assign  _seach_blockx_28_p_reset = p_reset;
   assign  _seach_blockx_28_m_clock = m_clock;
   assign  _seach_blockx_27_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in46:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_27_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00101110:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_27_in_do)
  begin
#1 if (_seach_blockx_27_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_27_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 41 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_27_in_do = (in_do|_reg_1);
   assign  _seach_blockx_27_p_reset = p_reset;
   assign  _seach_blockx_27_m_clock = m_clock;
   assign  _seach_blockx_26_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in45:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_26_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00101101:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_26_in_do)
  begin
#1 if (_seach_blockx_26_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_26_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 40 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_26_in_do = (in_do|_reg_1);
   assign  _seach_blockx_26_p_reset = p_reset;
   assign  _seach_blockx_26_m_clock = m_clock;
   assign  _seach_blockx_25_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in44:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_25_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00101100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_25_in_do)
  begin
#1 if (_seach_blockx_25_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_25_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 39 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_25_in_do = (in_do|_reg_1);
   assign  _seach_blockx_25_p_reset = p_reset;
   assign  _seach_blockx_25_m_clock = m_clock;
   assign  _seach_blockx_24_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in43:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_24_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00101011:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_24_in_do)
  begin
#1 if (_seach_blockx_24_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_24_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 38 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_24_in_do = (in_do|_reg_1);
   assign  _seach_blockx_24_p_reset = p_reset;
   assign  _seach_blockx_24_m_clock = m_clock;
   assign  _seach_blockx_23_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in42:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_23_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00101010:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_23_in_do)
  begin
#1 if (_seach_blockx_23_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_23_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 37 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_23_in_do = (in_do|_reg_1);
   assign  _seach_blockx_23_p_reset = p_reset;
   assign  _seach_blockx_23_m_clock = m_clock;
   assign  _seach_blockx_22_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in41:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_22_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00101001:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_22_in_do)
  begin
#1 if (_seach_blockx_22_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_22_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 36 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_22_in_do = (in_do|_reg_1);
   assign  _seach_blockx_22_p_reset = p_reset;
   assign  _seach_blockx_22_m_clock = m_clock;
   assign  _seach_blockx_21_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in40:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_21_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00101000:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_21_in_do)
  begin
#1 if (_seach_blockx_21_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_21_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 35 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_21_in_do = (in_do|_reg_1);
   assign  _seach_blockx_21_p_reset = p_reset;
   assign  _seach_blockx_21_m_clock = m_clock;
   assign  _seach_blockx_20_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in39:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_20_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00100111:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_20_in_do)
  begin
#1 if (_seach_blockx_20_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_20_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 34 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_20_in_do = (in_do|_reg_1);
   assign  _seach_blockx_20_p_reset = p_reset;
   assign  _seach_blockx_20_m_clock = m_clock;
   assign  _seach_blockx_19_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in38:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_19_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00100110:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_19_in_do)
  begin
#1 if (_seach_blockx_19_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_19_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 33 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_19_in_do = (in_do|_reg_1);
   assign  _seach_blockx_19_p_reset = p_reset;
   assign  _seach_blockx_19_m_clock = m_clock;
   assign  _seach_blockx_18_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in37:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_18_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00100101:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_18_in_do)
  begin
#1 if (_seach_blockx_18_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_18_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 32 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_18_in_do = (in_do|_reg_1);
   assign  _seach_blockx_18_p_reset = p_reset;
   assign  _seach_blockx_18_m_clock = m_clock;
   assign  _seach_blockx_17_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in36:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_17_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00100100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_17_in_do)
  begin
#1 if (_seach_blockx_17_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_17_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 31 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_17_in_do = (in_do|_reg_1);
   assign  _seach_blockx_17_p_reset = p_reset;
   assign  _seach_blockx_17_m_clock = m_clock;
   assign  _seach_blockx_16_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in35:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_16_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00100011:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_16_in_do)
  begin
#1 if (_seach_blockx_16_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_16_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 30 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_16_in_do = (in_do|_reg_1);
   assign  _seach_blockx_16_p_reset = p_reset;
   assign  _seach_blockx_16_m_clock = m_clock;
   assign  _seach_blockx_15_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in34:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_15_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00100010:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_15_in_do)
  begin
#1 if (_seach_blockx_15_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_15_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 29 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_15_in_do = (in_do|_reg_1);
   assign  _seach_blockx_15_p_reset = p_reset;
   assign  _seach_blockx_15_m_clock = m_clock;
   assign  _seach_blockx_14_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in33:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_14_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00100001:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_14_in_do)
  begin
#1 if (_seach_blockx_14_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_14_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 28 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_14_in_do = (in_do|_reg_1);
   assign  _seach_blockx_14_p_reset = p_reset;
   assign  _seach_blockx_14_m_clock = m_clock;
   assign  _seach_blockx_13_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in30:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_13_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00011110:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_13_in_do)
  begin
#1 if (_seach_blockx_13_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_13_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 27 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_13_in_do = (in_do|_reg_1);
   assign  _seach_blockx_13_p_reset = p_reset;
   assign  _seach_blockx_13_m_clock = m_clock;
   assign  _seach_blockx_12_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in29:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_12_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00011101:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_12_in_do)
  begin
#1 if (_seach_blockx_12_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_12_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 26 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_12_in_do = (in_do|_reg_1);
   assign  _seach_blockx_12_p_reset = p_reset;
   assign  _seach_blockx_12_m_clock = m_clock;
   assign  _seach_blockx_11_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in28:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_11_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00011100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_11_in_do)
  begin
#1 if (_seach_blockx_11_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_11_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 25 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_11_in_do = (in_do|_reg_1);
   assign  _seach_blockx_11_p_reset = p_reset;
   assign  _seach_blockx_11_m_clock = m_clock;
   assign  _seach_blockx_10_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in27:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_10_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00011011:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_10_in_do)
  begin
#1 if (_seach_blockx_10_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_10_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 24 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_10_in_do = (in_do|_reg_1);
   assign  _seach_blockx_10_p_reset = p_reset;
   assign  _seach_blockx_10_m_clock = m_clock;
   assign  _seach_blockx_9_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in26:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_9_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00011010:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_9_in_do)
  begin
#1 if (_seach_blockx_9_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_9_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 23 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_9_in_do = (in_do|_reg_1);
   assign  _seach_blockx_9_p_reset = p_reset;
   assign  _seach_blockx_9_m_clock = m_clock;
   assign  _seach_blockx_8_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in25:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_8_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00011001:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_8_in_do)
  begin
#1 if (_seach_blockx_8_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_8_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 22 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_8_in_do = (in_do|_reg_1);
   assign  _seach_blockx_8_p_reset = p_reset;
   assign  _seach_blockx_8_m_clock = m_clock;
   assign  _seach_blockx_7_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in24:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_7_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00011000:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_7_in_do)
  begin
#1 if (_seach_blockx_7_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_7_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 21 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_7_in_do = (in_do|_reg_1);
   assign  _seach_blockx_7_p_reset = p_reset;
   assign  _seach_blockx_7_m_clock = m_clock;
   assign  _seach_blockx_6_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in23:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_6_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00010111:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_6_in_do)
  begin
#1 if (_seach_blockx_6_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_6_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 20 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_6_in_do = (in_do|_reg_1);
   assign  _seach_blockx_6_p_reset = p_reset;
   assign  _seach_blockx_6_m_clock = m_clock;
   assign  _seach_blockx_5_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in22:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_5_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00010110:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_5_in_do)
  begin
#1 if (_seach_blockx_5_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_5_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 19 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_5_in_do = (in_do|_reg_1);
   assign  _seach_blockx_5_p_reset = p_reset;
   assign  _seach_blockx_5_m_clock = m_clock;
   assign  _seach_blockx_4_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in21:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_4_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00010101:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_4_in_do)
  begin
#1 if (_seach_blockx_4_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_4_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 18 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_4_in_do = (in_do|_reg_1);
   assign  _seach_blockx_4_p_reset = p_reset;
   assign  _seach_blockx_4_m_clock = m_clock;
   assign  _seach_blockx_3_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in20:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_3_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00010100:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_3_in_do)
  begin
#1 if (_seach_blockx_3_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_3_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 17 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_3_in_do = (in_do|_reg_1);
   assign  _seach_blockx_3_p_reset = p_reset;
   assign  _seach_blockx_3_m_clock = m_clock;
   assign  _seach_blockx_2_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in19:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_2_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00010011:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_2_in_do)
  begin
#1 if (_seach_blockx_2_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_2_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 16 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_2_in_do = (in_do|_reg_1);
   assign  _seach_blockx_2_p_reset = p_reset;
   assign  _seach_blockx_2_m_clock = m_clock;
   assign  _seach_blockx_1_map_block = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?data_in18:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;
   assign  _seach_blockx_1_now = 
// synthesis translate_off
// synopsys translate_off
((in_do|_reg_1))? 
// synthesis translate_on
// synopsys translate_on
(((in_do|_reg_1))?8'b00010010:8'b0)
// synthesis translate_off
// synopsys translate_off
:8'bx
// synthesis translate_on
// synopsys translate_on
;

// synthesis translate_off
// synopsys translate_off
always @(posedge _seach_blockx_1_in_do)
  begin
#1 if (_seach_blockx_1_in_do===1'bx)
 begin
$display("Warning: control hazard(seach:_seach_blockx_1_in_do) at %d",$time);
 end
#1 if ((((in_do|_reg_1))===1'bx) || (1'b1)===1'bx) $display("hazard ((in_do|_reg_1) || 1'b1) line 15 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  _seach_blockx_1_in_do = (in_do|_reg_1);
   assign  _seach_blockx_1_p_reset = p_reset;
   assign  _seach_blockx_1_m_clock = m_clock;
   assign  data_out17 = _seach_blockx_data_out;
   assign  data_out18 = _seach_blockx_1_data_out;
   assign  data_out19 = _seach_blockx_2_data_out;
   assign  data_out20 = _seach_blockx_3_data_out;
   assign  data_out21 = _seach_blockx_4_data_out;
   assign  data_out22 = _seach_blockx_5_data_out;
   assign  data_out23 = _seach_blockx_6_data_out;
   assign  data_out24 = _seach_blockx_7_data_out;
   assign  data_out25 = _seach_blockx_8_data_out;
   assign  data_out26 = _seach_blockx_9_data_out;
   assign  data_out27 = _seach_blockx_10_data_out;
   assign  data_out28 = _seach_blockx_11_data_out;
   assign  data_out29 = _seach_blockx_12_data_out;
   assign  data_out30 = _seach_blockx_13_data_out;
   assign  data_out33 = _seach_blockx_14_data_out;
   assign  data_out34 = _seach_blockx_15_data_out;
   assign  data_out35 = _seach_blockx_16_data_out;
   assign  data_out36 = _seach_blockx_17_data_out;
   assign  data_out37 = _seach_blockx_18_data_out;
   assign  data_out38 = _seach_blockx_19_data_out;
   assign  data_out39 = _seach_blockx_20_data_out;
   assign  data_out40 = _seach_blockx_21_data_out;
   assign  data_out41 = _seach_blockx_22_data_out;
   assign  data_out42 = _seach_blockx_23_data_out;
   assign  data_out43 = _seach_blockx_24_data_out;
   assign  data_out44 = _seach_blockx_25_data_out;
   assign  data_out45 = _seach_blockx_26_data_out;
   assign  data_out46 = _seach_blockx_27_data_out;
   assign  data_out49 = _seach_blockx_28_data_out;
   assign  data_out50 = _seach_blockx_29_data_out;
   assign  data_out51 = _seach_blockx_30_data_out;
   assign  data_out52 = _seach_blockx_31_data_out;
   assign  data_out53 = _seach_blockx_32_data_out;
   assign  data_out54 = _seach_blockx_33_data_out;
   assign  data_out55 = _seach_blockx_34_data_out;
   assign  data_out56 = _seach_blockx_35_data_out;
   assign  data_out57 = _seach_blockx_36_data_out;
   assign  data_out58 = _seach_blockx_37_data_out;
   assign  data_out59 = _seach_blockx_38_data_out;
   assign  data_out60 = _seach_blockx_39_data_out;
   assign  data_out61 = _seach_blockx_40_data_out;
   assign  data_out62 = _seach_blockx_41_data_out;
   assign  data_out65 = _seach_blockx_42_data_out;
   assign  data_out66 = _seach_blockx_43_data_out;
   assign  data_out67 = _seach_blockx_44_data_out;
   assign  data_out68 = _seach_blockx_45_data_out;
   assign  data_out69 = _seach_blockx_46_data_out;
   assign  data_out70 = _seach_blockx_47_data_out;
   assign  data_out71 = _seach_blockx_48_data_out;
   assign  data_out72 = _seach_blockx_49_data_out;
   assign  data_out73 = _seach_blockx_50_data_out;
   assign  data_out74 = _seach_blockx_51_data_out;
   assign  data_out75 = _seach_blockx_52_data_out;
   assign  data_out76 = _seach_blockx_53_data_out;
   assign  data_out77 = _seach_blockx_54_data_out;
   assign  data_out78 = _seach_blockx_55_data_out;
   assign  data_out81 = _seach_blockx_56_data_out;
   assign  data_out82 = _seach_blockx_57_data_out;
   assign  data_out83 = _seach_blockx_58_data_out;
   assign  data_out84 = _seach_blockx_59_data_out;
   assign  data_out85 = _seach_blockx_60_data_out;
   assign  data_out86 = _seach_blockx_61_data_out;
   assign  data_out87 = _seach_blockx_62_data_out;
   assign  data_out88 = _seach_blockx_63_data_out;
   assign  data_out89 = _seach_blockx_64_data_out;
   assign  data_out90 = _seach_blockx_65_data_out;
   assign  data_out91 = _seach_blockx_66_data_out;
   assign  data_out92 = _seach_blockx_67_data_out;
   assign  data_out93 = _seach_blockx_68_data_out;
   assign  data_out94 = _seach_blockx_69_data_out;
   assign  data_out97 = _seach_blockx_70_data_out;
   assign  data_out98 = _seach_blockx_71_data_out;
   assign  data_out99 = _seach_blockx_72_data_out;
   assign  data_out100 = _seach_blockx_73_data_out;
   assign  data_out101 = _seach_blockx_74_data_out;
   assign  data_out102 = _seach_blockx_75_data_out;
   assign  data_out103 = _seach_blockx_76_data_out;
   assign  data_out104 = _seach_blockx_77_data_out;
   assign  data_out105 = _seach_blockx_78_data_out;
   assign  data_out106 = _seach_blockx_79_data_out;
   assign  data_out107 = _seach_blockx_80_data_out;
   assign  data_out108 = _seach_blockx_81_data_out;
   assign  data_out109 = _seach_blockx_82_data_out;
   assign  data_out110 = _seach_blockx_83_data_out;
   assign  startplot = startplot_reg;
   assign  goalplot = goalplot_reg;

// synthesis translate_off
// synopsys translate_off
always @(posedge out_do)
  begin
#1 if (out_do===1'bx)
 begin
$display("Warning: control hazard(seach:out_do) at %d",$time);
 end
#1 if (((_reg_0)===1'bx) || (1'b1)===1'bx) $display("hazard (_reg_0 || 1'b1) line 104 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  out_do = _reg_0;

// synthesis translate_off
// synopsys translate_off
always @(posedge out_data)
  begin
#1 if (out_data===1'bx)
 begin
$display("Warning: control hazard(seach:out_data) at %d",$time);
 end
#1 if (((1'b1)===1'bx) || (1'b1)===1'bx) $display("hazard (1'b1 || 1'b1) line 8 at %d\n",$time);
 end

// synthesis translate_on
// synopsys translate_on
   assign  out_data = 1'b1;
always @(posedge m_clock or posedge p_reset)
  begin
if (p_reset)
     startplot_reg <= 8'b00000000;
else if ((in_do|_reg_1))
      startplot_reg <= (((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_seach_blockx_start|_seach_blockx_1_start)|_seach_blockx_2_start)|_seach_blockx_3_start)|_seach_blockx_4_start)|_seach_blockx_5_start)|_seach_blockx_6_start)|_seach_blockx_7_start)|_seach_blockx_8_start)|_seach_blockx_9_start)|_seach_blockx_10_start)|_seach_blockx_11_start)|_seach_blockx_12_start)|_seach_blockx_13_start)|_seach_blockx_14_start)|_seach_blockx_15_start)|_seach_blockx_16_start)|_seach_blockx_17_start)|_seach_blockx_18_start)|_seach_blockx_19_start)|_seach_blockx_20_start)|_seach_blockx_21_start)|_seach_blockx_22_start)|_seach_blockx_23_start)|_seach_blockx_24_start)|_seach_blockx_25_start)|_seach_blockx_26_start)|_seach_blockx_27_start)|_seach_blockx_28_start)|_seach_blockx_29_start)|_seach_blockx_30_start)|_seach_blockx_31_start)|_seach_blockx_32_start)|_seach_blockx_33_start)|_seach_blockx_34_start)|_seach_blockx_35_start)|_seach_blockx_36_start)|_seach_blockx_37_start)|_seach_blockx_38_start)|_seach_blockx_39_start)|_seach_blockx_40_start)|_seach_blockx_41_start)|_seach_blockx_42_start)|_seach_blockx_43_start)|_seach_blockx_44_start)|_seach_blockx_45_start)|_seach_blockx_46_start)|_seach_blockx_47_start)|_seach_blockx_48_start)|_seach_blockx_49_start)|_seach_blockx_50_start)|_seach_blockx_51_start)|_seach_blockx_52_start)|_seach_blockx_53_start)|_seach_blockx_54_start)|_seach_blockx_55_start)|_seach_blockx_56_start)|_seach_blockx_57_start)|_seach_blockx_58_start)|_seach_blockx_59_start)|_seach_blockx_60_start)|_seach_blockx_61_start)|_seach_blockx_62_start)|_seach_blockx_63_start)|_seach_blockx_64_start)|_seach_blockx_65_start)|_seach_blockx_66_start)|_seach_blockx_67_start)|_seach_blockx_68_start)|_seach_blockx_69_start)|_seach_blockx_70_start)|_seach_blockx_71_start)|_seach_blockx_72_start)|_seach_blockx_73_start)|_seach_blockx_74_start)|_seach_blockx_75_start)|_seach_blockx_76_start)|_seach_blockx_77_start)|_seach_blockx_78_start)|_seach_blockx_79_start)|_seach_blockx_80_start)|_seach_blockx_81_start)|_seach_blockx_82_start)|_seach_blockx_83_start);
end
always @(posedge m_clock or posedge p_reset)
  begin
if (p_reset)
     goalplot_reg <= 8'b00000000;
else if ((in_do|_reg_1))
      goalplot_reg <= (((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((((_seach_blockx_goal|_seach_blockx_1_goal)|_seach_blockx_2_goal)|_seach_blockx_3_goal)|_seach_blockx_4_goal)|_seach_blockx_5_goal)|_seach_blockx_6_goal)|_seach_blockx_7_goal)|_seach_blockx_8_goal)|_seach_blockx_9_goal)|_seach_blockx_10_goal)|_seach_blockx_11_goal)|_seach_blockx_12_goal)|_seach_blockx_13_goal)|_seach_blockx_14_goal)|_seach_blockx_15_goal)|_seach_blockx_16_goal)|_seach_blockx_17_goal)|_seach_blockx_18_goal)|_seach_blockx_19_goal)|_seach_blockx_20_goal)|_seach_blockx_21_goal)|_seach_blockx_22_goal)|_seach_blockx_23_goal)|_seach_blockx_24_goal)|_seach_blockx_25_goal)|_seach_blockx_26_goal)|_seach_blockx_27_goal)|_seach_blockx_28_goal)|_seach_blockx_29_goal)|_seach_blockx_30_goal)|_seach_blockx_31_goal)|_seach_blockx_32_goal)|_seach_blockx_33_goal)|_seach_blockx_34_goal)|_seach_blockx_35_goal)|_seach_blockx_36_goal)|_seach_blockx_37_goal)|_seach_blockx_38_goal)|_seach_blockx_39_goal)|_seach_blockx_40_goal)|_seach_blockx_41_goal)|_seach_blockx_42_goal)|_seach_blockx_43_goal)|_seach_blockx_44_goal)|_seach_blockx_45_goal)|_seach_blockx_46_goal)|_seach_blockx_47_goal)|_seach_blockx_48_goal)|_seach_blockx_49_goal)|_seach_blockx_50_goal)|_seach_blockx_51_goal)|_seach_blockx_52_goal)|_seach_blockx_53_goal)|_seach_blockx_54_goal)|_seach_blockx_55_goal)|_seach_blockx_56_goal)|_seach_blockx_57_goal)|_seach_blockx_58_goal)|_seach_blockx_59_goal)|_seach_blockx_60_goal)|_seach_blockx_61_goal)|_seach_blockx_62_goal)|_seach_blockx_63_goal)|_seach_blockx_64_goal)|_seach_blockx_65_goal)|_seach_blockx_66_goal)|_seach_blockx_67_goal)|_seach_blockx_68_goal)|_seach_blockx_69_goal)|_seach_blockx_70_goal)|_seach_blockx_71_goal)|_seach_blockx_72_goal)|_seach_blockx_73_goal)|_seach_blockx_74_goal)|_seach_blockx_75_goal)|_seach_blockx_76_goal)|_seach_blockx_77_goal)|_seach_blockx_78_goal)|_seach_blockx_79_goal)|_seach_blockx_80_goal)|_seach_blockx_81_goal)|_seach_blockx_82_goal)|_seach_blockx_83_goal);
end
always @(posedge m_clock or posedge p_reset)
  begin
if (p_reset)
     _reg_0 <= 1'b0;
else if ((in_do|(_reg_0|_reg_1)))
      _reg_0 <= (_reg_1|in_do);
end
always @(posedge m_clock or posedge p_reset)
  begin
if (p_reset)
     _reg_1 <= 1'b0;
else if (_reg_1)
      _reg_1 <= 1'b0;
end
endmodule

/*Produced by NSL Core(version=20240424), IP ARCH, Inc. Tue May 21 04:56:16 2024
 Licensed to :EVALUATION USER*/
